module rom_num2(clock, address, q);     // ROM-stored RGB bitmap for "2"
input clock;
output [7:0] q;
input [10:0] address;
reg [7:0] dout;
reg [7:0] ram [2047:0];
assign q = dout;

initial begin
  ram[0]  = 255;
  ram[1]  = 255;
  ram[2]  = 255;
  ram[3]  = 255;
  ram[4]  = 255;
  ram[5]  = 255;
  ram[6]  = 255;
  ram[7]  = 255;
  ram[8]  = 255;
  ram[9]  = 255;
  ram[10]  = 255;
  ram[11]  = 255;
  ram[12]  = 255;
  ram[13]  = 255;
  ram[14]  = 255;
  ram[15]  = 255;
  ram[16]  = 255;
  ram[17]  = 255;
  ram[18]  = 255;
  ram[19]  = 255;
  ram[20]  = 255;
  ram[21]  = 255;
  ram[22]  = 255;
  ram[23]  = 255;
  ram[24]  = 255;
  ram[25]  = 255;
  ram[26]  = 255;
  ram[27]  = 255;
  ram[28]  = 255;
  ram[29]  = 255;
  ram[30]  = 255;
  ram[31]  = 255;
  ram[32]  = 255;
  ram[33]  = 255;
  ram[34]  = 255;
  ram[35]  = 255;
  ram[36]  = 255;
  ram[37]  = 255;
  ram[38]  = 255;
  ram[39]  = 255;
  ram[40]  = 255;
  ram[41]  = 255;
  ram[42]  = 255;
  ram[43]  = 255;
  ram[44]  = 255;
  ram[45]  = 255;
  ram[46]  = 255;
  ram[47]  = 255;
  ram[48]  = 255;
  ram[49]  = 255;
  ram[50]  = 255;
  ram[51]  = 255;
  ram[52]  = 255;
  ram[53]  = 255;
  ram[54]  = 255;
  ram[55]  = 255;
  ram[56]  = 255;
  ram[57]  = 255;
  ram[58]  = 255;
  ram[59]  = 255;
  ram[60]  = 255;
  ram[61]  = 255;
  ram[62]  = 255;
  ram[63]  = 255;
  ram[64]  = 255;
  ram[65]  = 255;
  ram[66]  = 255;
  ram[67]  = 255;
  ram[68]  = 255;
  ram[69]  = 255;
  ram[70]  = 255;
  ram[71]  = 255;
  ram[72]  = 255;
  ram[73]  = 255;
  ram[74]  = 255;
  ram[75]  = 255;
  ram[76]  = 255;
  ram[77]  = 255;
  ram[78]  = 255;
  ram[79]  = 255;
  ram[80]  = 255;
  ram[81]  = 255;
  ram[82]  = 255;
  ram[83]  = 255;
  ram[84]  = 255;
  ram[85]  = 255;
  ram[86]  = 255;
  ram[87]  = 255;
  ram[88]  = 255;
  ram[89]  = 255;
  ram[90]  = 255;
  ram[91]  = 255;
  ram[92]  = 255;
  ram[93]  = 255;
  ram[94]  = 255;
  ram[95]  = 255;
  ram[96]  = 255;
  ram[97]  = 255;
  ram[98]  = 255;
  ram[99]  = 255;
  ram[100]  = 255;
  ram[101]  = 255;
  ram[102]  = 255;
  ram[103]  = 255;
  ram[104]  = 255;
  ram[105]  = 255;
  ram[106]  = 255;
  ram[107]  = 255;
  ram[108]  = 255;
  ram[109]  = 255;
  ram[110]  = 255;
  ram[111]  = 255;
  ram[112]  = 255;
  ram[113]  = 255;
  ram[114]  = 255;
  ram[115]  = 255;
  ram[116]  = 255;
  ram[117]  = 255;
  ram[118]  = 255;
  ram[119]  = 255;
  ram[120]  = 255;
  ram[121]  = 255;
  ram[122]  = 255;
  ram[123]  = 255;
  ram[124]  = 255;
  ram[125]  = 255;
  ram[126]  = 255;
  ram[127]  = 255;
  ram[128]  = 255;
  ram[129]  = 255;
  ram[130]  = 255;
  ram[131]  = 255;
  ram[132]  = 255;
  ram[133]  = 255;
  ram[134]  = 255;
  ram[135]  = 255;
  ram[136]  = 255;
  ram[137]  = 255;
  ram[138]  = 255;
  ram[139]  = 255;
  ram[140]  = 255;
  ram[141]  = 255;
  ram[142]  = 255;
  ram[143]  = 255;
  ram[144]  = 255;
  ram[145]  = 255;
  ram[146]  = 255;
  ram[147]  = 255;
  ram[148]  = 255;
  ram[149]  = 255;
  ram[150]  = 255;
  ram[151]  = 255;
  ram[152]  = 255;
  ram[153]  = 255;
  ram[154]  = 255;
  ram[155]  = 255;
  ram[156]  = 255;
  ram[157]  = 255;
  ram[158]  = 255;
  ram[159]  = 255;
  ram[160]  = 255;
  ram[161]  = 255;
  ram[162]  = 255;
  ram[163]  = 255;
  ram[164]  = 255;
  ram[165]  = 255;
  ram[166]  = 255;
  ram[167]  = 255;
  ram[168]  = 255;
  ram[169]  = 255;
  ram[170]  = 255;
  ram[171]  = 255;
  ram[172]  = 255;
  ram[173]  = 255;
  ram[174]  = 255;
  ram[175]  = 255;
  ram[176]  = 255;
  ram[177]  = 255;
  ram[178]  = 255;
  ram[179]  = 255;
  ram[180]  = 255;
  ram[181]  = 255;
  ram[182]  = 255;
  ram[183]  = 255;
  ram[184]  = 255;
  ram[185]  = 255;
  ram[186]  = 255;
  ram[187]  = 255;
  ram[188]  = 255;
  ram[189]  = 255;
  ram[190]  = 255;
  ram[191]  = 255;
  ram[192]  = 255;
  ram[193]  = 255;
  ram[194]  = 255;
  ram[195]  = 255;
  ram[196]  = 255;
  ram[197]  = 255;
  ram[198]  = 255;
  ram[199]  = 255;
  ram[200]  = 255;
  ram[201]  = 255;
  ram[202]  = 255;
  ram[203]  = 255;
  ram[204]  = 255;
  ram[205]  = 255;
  ram[206]  = 255;
  ram[207]  = 255;
  ram[208]  = 255;
  ram[209]  = 255;
  ram[210]  = 255;
  ram[211]  = 255;
  ram[212]  = 255;
  ram[213]  = 255;
  ram[214]  = 255;
  ram[215]  = 255;
  ram[216]  = 255;
  ram[217]  = 255;
  ram[218]  = 255;
  ram[219]  = 255;
  ram[220]  = 255;
  ram[221]  = 255;
  ram[222]  = 255;
  ram[223]  = 255;
  ram[224]  = 255;
  ram[225]  = 255;
  ram[226]  = 255;
  ram[227]  = 255;
  ram[228]  = 255;
  ram[229]  = 255;
  ram[230]  = 255;
  ram[231]  = 255;
  ram[232]  = 255;
  ram[233]  = 255;
  ram[234]  = 255;
  ram[235]  = 255;
  ram[236]  = 255;
  ram[237]  = 255;
  ram[238]  = 255;
  ram[239]  = 255;
  ram[240]  = 255;
  ram[241]  = 255;
  ram[242]  = 255;
  ram[243]  = 255;
  ram[244]  = 255;
  ram[245]  = 255;
  ram[246]  = 255;
  ram[247]  = 255;
  ram[248]  = 255;
  ram[249]  = 255;
  ram[250]  = 255;
  ram[251]  = 255;
  ram[252]  = 255;
  ram[253]  = 255;
  ram[254]  = 255;
  ram[255]  = 255;
  ram[256]  = 255;
  ram[257]  = 255;
  ram[258]  = 255;
  ram[259]  = 255;
  ram[260]  = 255;
  ram[261]  = 255;
  ram[262]  = 255;
  ram[263]  = 255;
  ram[264]  = 255;
  ram[265]  = 255;
  ram[266]  = 255;
  ram[267]  = 255;
  ram[268]  = 255;
  ram[269]  = 255;
  ram[270]  = 255;
  ram[271]  = 255;
  ram[272]  = 255;
  ram[273]  = 255;
  ram[274]  = 255;
  ram[275]  = 255;
  ram[276]  = 255;
  ram[277]  = 255;
  ram[278]  = 255;
  ram[279]  = 255;
  ram[280]  = 255;
  ram[281]  = 255;
  ram[282]  = 255;
  ram[283]  = 255;
  ram[284]  = 255;
  ram[285]  = 255;
  ram[286]  = 255;
  ram[287]  = 255;
  ram[288]  = 255;
  ram[289]  = 255;
  ram[290]  = 255;
  ram[291]  = 255;
  ram[292]  = 255;
  ram[293]  = 255;
  ram[294]  = 255;
  ram[295]  = 255;
  ram[296]  = 255;
  ram[297]  = 255;
  ram[298]  = 255;
  ram[299]  = 255;
  ram[300]  = 255;
  ram[301]  = 255;
  ram[302]  = 255;
  ram[303]  = 255;
  ram[304]  = 255;
  ram[305]  = 255;
  ram[306]  = 255;
  ram[307]  = 255;
  ram[308]  = 255;
  ram[309]  = 255;
  ram[310]  = 255;
  ram[311]  = 255;
  ram[312]  = 255;
  ram[313]  = 255;
  ram[314]  = 255;
  ram[315]  = 255;
  ram[316]  = 255;
  ram[317]  = 255;
  ram[318]  = 255;
  ram[319]  = 255;
  ram[320]  = 255;
  ram[321]  = 255;
  ram[322]  = 255;
  ram[323]  = 255;
  ram[324]  = 255;
  ram[325]  = 255;
  ram[326]  = 255;
  ram[327]  = 255;
  ram[328]  = 255;
  ram[329]  = 255;
  ram[330]  = 255;
  ram[331]  = 255;
  ram[332]  = 255;
  ram[333]  = 255;
  ram[334]  = 255;
  ram[335]  = 221;
  ram[336]  = 137;
  ram[337]  = 71;
  ram[338]  = 71;
  ram[339]  = 71;
  ram[340]  = 122;
  ram[341]  = 195;
  ram[342]  = 255;
  ram[343]  = 255;
  ram[344]  = 255;
  ram[345]  = 255;
  ram[346]  = 255;
  ram[347]  = 255;
  ram[348]  = 255;
  ram[349]  = 255;
  ram[350]  = 255;
  ram[351]  = 255;
  ram[352]  = 255;
  ram[353]  = 255;
  ram[354]  = 255;
  ram[355]  = 255;
  ram[356]  = 255;
  ram[357]  = 255;
  ram[358]  = 255;
  ram[359]  = 255;
  ram[360]  = 255;
  ram[361]  = 255;
  ram[362]  = 255;
  ram[363]  = 255;
  ram[364]  = 255;
  ram[365]  = 255;
  ram[366]  = 255;
  ram[367]  = 255;
  ram[368]  = 255;
  ram[369]  = 255;
  ram[370]  = 255;
  ram[371]  = 255;
  ram[372]  = 255;
  ram[373]  = 255;
  ram[374]  = 122;
  ram[375]  = 0;
  ram[376]  = 0;
  ram[377]  = 0;
  ram[378]  = 0;
  ram[379]  = 0;
  ram[380]  = 0;
  ram[381]  = 0;
  ram[382]  = 71;
  ram[383]  = 236;
  ram[384]  = 255;
  ram[385]  = 255;
  ram[386]  = 255;
  ram[387]  = 255;
  ram[388]  = 255;
  ram[389]  = 255;
  ram[390]  = 255;
  ram[391]  = 255;
  ram[392]  = 255;
  ram[393]  = 255;
  ram[394]  = 255;
  ram[395]  = 255;
  ram[396]  = 255;
  ram[397]  = 255;
  ram[398]  = 255;
  ram[399]  = 255;
  ram[400]  = 255;
  ram[401]  = 255;
  ram[402]  = 255;
  ram[403]  = 255;
  ram[404]  = 255;
  ram[405]  = 255;
  ram[406]  = 255;
  ram[407]  = 255;
  ram[408]  = 255;
  ram[409]  = 255;
  ram[410]  = 255;
  ram[411]  = 255;
  ram[412]  = 255;
  ram[413]  = 152;
  ram[414]  = 0;
  ram[415]  = 0;
  ram[416]  = 71;
  ram[417]  = 137;
  ram[418]  = 137;
  ram[419]  = 137;
  ram[420]  = 35;
  ram[421]  = 0;
  ram[422]  = 0;
  ram[423]  = 52;
  ram[424]  = 255;
  ram[425]  = 255;
  ram[426]  = 255;
  ram[427]  = 255;
  ram[428]  = 255;
  ram[429]  = 255;
  ram[430]  = 255;
  ram[431]  = 255;
  ram[432]  = 255;
  ram[433]  = 255;
  ram[434]  = 255;
  ram[435]  = 255;
  ram[436]  = 255;
  ram[437]  = 255;
  ram[438]  = 255;
  ram[439]  = 255;
  ram[440]  = 255;
  ram[441]  = 255;
  ram[442]  = 255;
  ram[443]  = 255;
  ram[444]  = 255;
  ram[445]  = 255;
  ram[446]  = 255;
  ram[447]  = 255;
  ram[448]  = 255;
  ram[449]  = 255;
  ram[450]  = 255;
  ram[451]  = 255;
  ram[452]  = 255;
  ram[453]  = 137;
  ram[454]  = 52;
  ram[455]  = 195;
  ram[456]  = 255;
  ram[457]  = 255;
  ram[458]  = 255;
  ram[459]  = 255;
  ram[460]  = 255;
  ram[461]  = 105;
  ram[462]  = 0;
  ram[463]  = 0;
  ram[464]  = 167;
  ram[465]  = 255;
  ram[466]  = 255;
  ram[467]  = 255;
  ram[468]  = 255;
  ram[469]  = 255;
  ram[470]  = 255;
  ram[471]  = 255;
  ram[472]  = 255;
  ram[473]  = 255;
  ram[474]  = 255;
  ram[475]  = 255;
  ram[476]  = 255;
  ram[477]  = 255;
  ram[478]  = 255;
  ram[479]  = 255;
  ram[480]  = 255;
  ram[481]  = 255;
  ram[482]  = 255;
  ram[483]  = 255;
  ram[484]  = 255;
  ram[485]  = 255;
  ram[486]  = 255;
  ram[487]  = 255;
  ram[488]  = 255;
  ram[489]  = 255;
  ram[490]  = 255;
  ram[491]  = 255;
  ram[492]  = 255;
  ram[493]  = 181;
  ram[494]  = 236;
  ram[495]  = 255;
  ram[496]  = 255;
  ram[497]  = 255;
  ram[498]  = 255;
  ram[499]  = 255;
  ram[500]  = 255;
  ram[501]  = 236;
  ram[502]  = 0;
  ram[503]  = 0;
  ram[504]  = 87;
  ram[505]  = 255;
  ram[506]  = 255;
  ram[507]  = 255;
  ram[508]  = 255;
  ram[509]  = 255;
  ram[510]  = 255;
  ram[511]  = 255;
  ram[512]  = 255;
  ram[513]  = 255;
  ram[514]  = 255;
  ram[515]  = 255;
  ram[516]  = 255;
  ram[517]  = 255;
  ram[518]  = 255;
  ram[519]  = 255;
  ram[520]  = 255;
  ram[521]  = 255;
  ram[522]  = 255;
  ram[523]  = 255;
  ram[524]  = 255;
  ram[525]  = 255;
  ram[526]  = 255;
  ram[527]  = 255;
  ram[528]  = 255;
  ram[529]  = 255;
  ram[530]  = 255;
  ram[531]  = 255;
  ram[532]  = 255;
  ram[533]  = 255;
  ram[534]  = 255;
  ram[535]  = 255;
  ram[536]  = 255;
  ram[537]  = 255;
  ram[538]  = 255;
  ram[539]  = 255;
  ram[540]  = 255;
  ram[541]  = 255;
  ram[542]  = 71;
  ram[543]  = 0;
  ram[544]  = 71;
  ram[545]  = 255;
  ram[546]  = 255;
  ram[547]  = 255;
  ram[548]  = 255;
  ram[549]  = 255;
  ram[550]  = 255;
  ram[551]  = 255;
  ram[552]  = 255;
  ram[553]  = 255;
  ram[554]  = 255;
  ram[555]  = 255;
  ram[556]  = 255;
  ram[557]  = 255;
  ram[558]  = 255;
  ram[559]  = 255;
  ram[560]  = 255;
  ram[561]  = 255;
  ram[562]  = 255;
  ram[563]  = 255;
  ram[564]  = 255;
  ram[565]  = 255;
  ram[566]  = 255;
  ram[567]  = 255;
  ram[568]  = 255;
  ram[569]  = 255;
  ram[570]  = 255;
  ram[571]  = 255;
  ram[572]  = 255;
  ram[573]  = 255;
  ram[574]  = 255;
  ram[575]  = 255;
  ram[576]  = 255;
  ram[577]  = 255;
  ram[578]  = 255;
  ram[579]  = 255;
  ram[580]  = 255;
  ram[581]  = 255;
  ram[582]  = 71;
  ram[583]  = 0;
  ram[584]  = 71;
  ram[585]  = 255;
  ram[586]  = 255;
  ram[587]  = 255;
  ram[588]  = 255;
  ram[589]  = 255;
  ram[590]  = 255;
  ram[591]  = 255;
  ram[592]  = 255;
  ram[593]  = 255;
  ram[594]  = 255;
  ram[595]  = 255;
  ram[596]  = 255;
  ram[597]  = 255;
  ram[598]  = 255;
  ram[599]  = 255;
  ram[600]  = 255;
  ram[601]  = 255;
  ram[602]  = 255;
  ram[603]  = 255;
  ram[604]  = 255;
  ram[605]  = 255;
  ram[606]  = 255;
  ram[607]  = 255;
  ram[608]  = 255;
  ram[609]  = 255;
  ram[610]  = 255;
  ram[611]  = 255;
  ram[612]  = 255;
  ram[613]  = 255;
  ram[614]  = 255;
  ram[615]  = 255;
  ram[616]  = 255;
  ram[617]  = 255;
  ram[618]  = 255;
  ram[619]  = 255;
  ram[620]  = 255;
  ram[621]  = 255;
  ram[622]  = 0;
  ram[623]  = 0;
  ram[624]  = 105;
  ram[625]  = 255;
  ram[626]  = 255;
  ram[627]  = 255;
  ram[628]  = 255;
  ram[629]  = 255;
  ram[630]  = 255;
  ram[631]  = 255;
  ram[632]  = 255;
  ram[633]  = 255;
  ram[634]  = 255;
  ram[635]  = 255;
  ram[636]  = 255;
  ram[637]  = 255;
  ram[638]  = 255;
  ram[639]  = 255;
  ram[640]  = 255;
  ram[641]  = 255;
  ram[642]  = 255;
  ram[643]  = 255;
  ram[644]  = 255;
  ram[645]  = 255;
  ram[646]  = 255;
  ram[647]  = 255;
  ram[648]  = 255;
  ram[649]  = 255;
  ram[650]  = 255;
  ram[651]  = 255;
  ram[652]  = 255;
  ram[653]  = 255;
  ram[654]  = 255;
  ram[655]  = 255;
  ram[656]  = 255;
  ram[657]  = 255;
  ram[658]  = 255;
  ram[659]  = 255;
  ram[660]  = 255;
  ram[661]  = 152;
  ram[662]  = 0;
  ram[663]  = 0;
  ram[664]  = 181;
  ram[665]  = 255;
  ram[666]  = 255;
  ram[667]  = 255;
  ram[668]  = 255;
  ram[669]  = 255;
  ram[670]  = 255;
  ram[671]  = 255;
  ram[672]  = 255;
  ram[673]  = 255;
  ram[674]  = 255;
  ram[675]  = 255;
  ram[676]  = 255;
  ram[677]  = 255;
  ram[678]  = 255;
  ram[679]  = 255;
  ram[680]  = 255;
  ram[681]  = 255;
  ram[682]  = 255;
  ram[683]  = 255;
  ram[684]  = 255;
  ram[685]  = 255;
  ram[686]  = 255;
  ram[687]  = 255;
  ram[688]  = 255;
  ram[689]  = 255;
  ram[690]  = 255;
  ram[691]  = 255;
  ram[692]  = 255;
  ram[693]  = 255;
  ram[694]  = 255;
  ram[695]  = 255;
  ram[696]  = 255;
  ram[697]  = 255;
  ram[698]  = 255;
  ram[699]  = 255;
  ram[700]  = 208;
  ram[701]  = 17;
  ram[702]  = 0;
  ram[703]  = 52;
  ram[704]  = 255;
  ram[705]  = 255;
  ram[706]  = 255;
  ram[707]  = 255;
  ram[708]  = 255;
  ram[709]  = 255;
  ram[710]  = 255;
  ram[711]  = 255;
  ram[712]  = 255;
  ram[713]  = 255;
  ram[714]  = 255;
  ram[715]  = 255;
  ram[716]  = 255;
  ram[717]  = 255;
  ram[718]  = 255;
  ram[719]  = 255;
  ram[720]  = 255;
  ram[721]  = 255;
  ram[722]  = 255;
  ram[723]  = 255;
  ram[724]  = 255;
  ram[725]  = 255;
  ram[726]  = 255;
  ram[727]  = 255;
  ram[728]  = 255;
  ram[729]  = 255;
  ram[730]  = 255;
  ram[731]  = 255;
  ram[732]  = 255;
  ram[733]  = 255;
  ram[734]  = 255;
  ram[735]  = 255;
  ram[736]  = 255;
  ram[737]  = 255;
  ram[738]  = 255;
  ram[739]  = 181;
  ram[740]  = 17;
  ram[741]  = 0;
  ram[742]  = 17;
  ram[743]  = 208;
  ram[744]  = 255;
  ram[745]  = 255;
  ram[746]  = 255;
  ram[747]  = 255;
  ram[748]  = 255;
  ram[749]  = 255;
  ram[750]  = 255;
  ram[751]  = 255;
  ram[752]  = 255;
  ram[753]  = 255;
  ram[754]  = 255;
  ram[755]  = 255;
  ram[756]  = 255;
  ram[757]  = 255;
  ram[758]  = 255;
  ram[759]  = 255;
  ram[760]  = 255;
  ram[761]  = 255;
  ram[762]  = 255;
  ram[763]  = 255;
  ram[764]  = 255;
  ram[765]  = 255;
  ram[766]  = 255;
  ram[767]  = 255;
  ram[768]  = 255;
  ram[769]  = 255;
  ram[770]  = 255;
  ram[771]  = 255;
  ram[772]  = 255;
  ram[773]  = 255;
  ram[774]  = 255;
  ram[775]  = 255;
  ram[776]  = 255;
  ram[777]  = 255;
  ram[778]  = 137;
  ram[779]  = 0;
  ram[780]  = 0;
  ram[781]  = 17;
  ram[782]  = 208;
  ram[783]  = 255;
  ram[784]  = 255;
  ram[785]  = 255;
  ram[786]  = 255;
  ram[787]  = 255;
  ram[788]  = 255;
  ram[789]  = 255;
  ram[790]  = 255;
  ram[791]  = 255;
  ram[792]  = 255;
  ram[793]  = 255;
  ram[794]  = 255;
  ram[795]  = 255;
  ram[796]  = 255;
  ram[797]  = 255;
  ram[798]  = 255;
  ram[799]  = 255;
  ram[800]  = 255;
  ram[801]  = 255;
  ram[802]  = 255;
  ram[803]  = 255;
  ram[804]  = 255;
  ram[805]  = 255;
  ram[806]  = 255;
  ram[807]  = 255;
  ram[808]  = 255;
  ram[809]  = 255;
  ram[810]  = 255;
  ram[811]  = 255;
  ram[812]  = 255;
  ram[813]  = 255;
  ram[814]  = 255;
  ram[815]  = 255;
  ram[816]  = 221;
  ram[817]  = 52;
  ram[818]  = 0;
  ram[819]  = 0;
  ram[820]  = 52;
  ram[821]  = 221;
  ram[822]  = 255;
  ram[823]  = 255;
  ram[824]  = 255;
  ram[825]  = 255;
  ram[826]  = 255;
  ram[827]  = 255;
  ram[828]  = 255;
  ram[829]  = 255;
  ram[830]  = 255;
  ram[831]  = 255;
  ram[832]  = 255;
  ram[833]  = 255;
  ram[834]  = 255;
  ram[835]  = 255;
  ram[836]  = 255;
  ram[837]  = 255;
  ram[838]  = 255;
  ram[839]  = 255;
  ram[840]  = 255;
  ram[841]  = 255;
  ram[842]  = 255;
  ram[843]  = 255;
  ram[844]  = 255;
  ram[845]  = 255;
  ram[846]  = 255;
  ram[847]  = 255;
  ram[848]  = 255;
  ram[849]  = 255;
  ram[850]  = 255;
  ram[851]  = 255;
  ram[852]  = 255;
  ram[853]  = 255;
  ram[854]  = 255;
  ram[855]  = 208;
  ram[856]  = 17;
  ram[857]  = 0;
  ram[858]  = 0;
  ram[859]  = 137;
  ram[860]  = 255;
  ram[861]  = 255;
  ram[862]  = 255;
  ram[863]  = 255;
  ram[864]  = 255;
  ram[865]  = 255;
  ram[866]  = 255;
  ram[867]  = 255;
  ram[868]  = 255;
  ram[869]  = 255;
  ram[870]  = 255;
  ram[871]  = 255;
  ram[872]  = 255;
  ram[873]  = 255;
  ram[874]  = 255;
  ram[875]  = 255;
  ram[876]  = 255;
  ram[877]  = 255;
  ram[878]  = 255;
  ram[879]  = 255;
  ram[880]  = 255;
  ram[881]  = 255;
  ram[882]  = 255;
  ram[883]  = 255;
  ram[884]  = 255;
  ram[885]  = 255;
  ram[886]  = 255;
  ram[887]  = 255;
  ram[888]  = 255;
  ram[889]  = 255;
  ram[890]  = 255;
  ram[891]  = 255;
  ram[892]  = 255;
  ram[893]  = 255;
  ram[894]  = 181;
  ram[895]  = 0;
  ram[896]  = 0;
  ram[897]  = 17;
  ram[898]  = 195;
  ram[899]  = 255;
  ram[900]  = 255;
  ram[901]  = 255;
  ram[902]  = 255;
  ram[903]  = 255;
  ram[904]  = 255;
  ram[905]  = 255;
  ram[906]  = 255;
  ram[907]  = 255;
  ram[908]  = 255;
  ram[909]  = 255;
  ram[910]  = 255;
  ram[911]  = 255;
  ram[912]  = 255;
  ram[913]  = 255;
  ram[914]  = 255;
  ram[915]  = 255;
  ram[916]  = 255;
  ram[917]  = 255;
  ram[918]  = 255;
  ram[919]  = 255;
  ram[920]  = 255;
  ram[921]  = 255;
  ram[922]  = 255;
  ram[923]  = 255;
  ram[924]  = 255;
  ram[925]  = 255;
  ram[926]  = 255;
  ram[927]  = 255;
  ram[928]  = 255;
  ram[929]  = 255;
  ram[930]  = 255;
  ram[931]  = 255;
  ram[932]  = 255;
  ram[933]  = 208;
  ram[934]  = 17;
  ram[935]  = 0;
  ram[936]  = 52;
  ram[937]  = 236;
  ram[938]  = 255;
  ram[939]  = 255;
  ram[940]  = 255;
  ram[941]  = 255;
  ram[942]  = 255;
  ram[943]  = 255;
  ram[944]  = 255;
  ram[945]  = 255;
  ram[946]  = 255;
  ram[947]  = 255;
  ram[948]  = 255;
  ram[949]  = 255;
  ram[950]  = 255;
  ram[951]  = 255;
  ram[952]  = 255;
  ram[953]  = 255;
  ram[954]  = 255;
  ram[955]  = 255;
  ram[956]  = 255;
  ram[957]  = 255;
  ram[958]  = 255;
  ram[959]  = 255;
  ram[960]  = 255;
  ram[961]  = 255;
  ram[962]  = 255;
  ram[963]  = 255;
  ram[964]  = 255;
  ram[965]  = 255;
  ram[966]  = 255;
  ram[967]  = 255;
  ram[968]  = 255;
  ram[969]  = 255;
  ram[970]  = 255;
  ram[971]  = 255;
  ram[972]  = 255;
  ram[973]  = 71;
  ram[974]  = 0;
  ram[975]  = 35;
  ram[976]  = 236;
  ram[977]  = 255;
  ram[978]  = 255;
  ram[979]  = 255;
  ram[980]  = 255;
  ram[981]  = 255;
  ram[982]  = 255;
  ram[983]  = 255;
  ram[984]  = 255;
  ram[985]  = 255;
  ram[986]  = 255;
  ram[987]  = 255;
  ram[988]  = 255;
  ram[989]  = 255;
  ram[990]  = 255;
  ram[991]  = 255;
  ram[992]  = 255;
  ram[993]  = 255;
  ram[994]  = 255;
  ram[995]  = 255;
  ram[996]  = 255;
  ram[997]  = 255;
  ram[998]  = 255;
  ram[999]  = 255;
  ram[1000]  = 255;
  ram[1001]  = 255;
  ram[1002]  = 255;
  ram[1003]  = 255;
  ram[1004]  = 255;
  ram[1005]  = 255;
  ram[1006]  = 255;
  ram[1007]  = 255;
  ram[1008]  = 255;
  ram[1009]  = 255;
  ram[1010]  = 255;
  ram[1011]  = 255;
  ram[1012]  = 221;
  ram[1013]  = 0;
  ram[1014]  = 0;
  ram[1015]  = 152;
  ram[1016]  = 255;
  ram[1017]  = 255;
  ram[1018]  = 255;
  ram[1019]  = 255;
  ram[1020]  = 255;
  ram[1021]  = 255;
  ram[1022]  = 255;
  ram[1023]  = 255;
  ram[1024]  = 255;
  ram[1025]  = 255;
  ram[1026]  = 255;
  ram[1027]  = 255;
  ram[1028]  = 255;
  ram[1029]  = 255;
  ram[1030]  = 255;
  ram[1031]  = 255;
  ram[1032]  = 255;
  ram[1033]  = 255;
  ram[1034]  = 255;
  ram[1035]  = 255;
  ram[1036]  = 255;
  ram[1037]  = 255;
  ram[1038]  = 255;
  ram[1039]  = 255;
  ram[1040]  = 255;
  ram[1041]  = 255;
  ram[1042]  = 255;
  ram[1043]  = 255;
  ram[1044]  = 255;
  ram[1045]  = 255;
  ram[1046]  = 255;
  ram[1047]  = 255;
  ram[1048]  = 255;
  ram[1049]  = 255;
  ram[1050]  = 255;
  ram[1051]  = 255;
  ram[1052]  = 181;
  ram[1053]  = 0;
  ram[1054]  = 0;
  ram[1055]  = 152;
  ram[1056]  = 195;
  ram[1057]  = 195;
  ram[1058]  = 195;
  ram[1059]  = 195;
  ram[1060]  = 195;
  ram[1061]  = 195;
  ram[1062]  = 195;
  ram[1063]  = 195;
  ram[1064]  = 195;
  ram[1065]  = 221;
  ram[1066]  = 255;
  ram[1067]  = 255;
  ram[1068]  = 255;
  ram[1069]  = 255;
  ram[1070]  = 255;
  ram[1071]  = 255;
  ram[1072]  = 255;
  ram[1073]  = 255;
  ram[1074]  = 255;
  ram[1075]  = 255;
  ram[1076]  = 255;
  ram[1077]  = 255;
  ram[1078]  = 255;
  ram[1079]  = 255;
  ram[1080]  = 255;
  ram[1081]  = 255;
  ram[1082]  = 255;
  ram[1083]  = 255;
  ram[1084]  = 255;
  ram[1085]  = 255;
  ram[1086]  = 255;
  ram[1087]  = 255;
  ram[1088]  = 255;
  ram[1089]  = 255;
  ram[1090]  = 255;
  ram[1091]  = 255;
  ram[1092]  = 137;
  ram[1093]  = 0;
  ram[1094]  = 0;
  ram[1095]  = 0;
  ram[1096]  = 0;
  ram[1097]  = 0;
  ram[1098]  = 0;
  ram[1099]  = 0;
  ram[1100]  = 0;
  ram[1101]  = 0;
  ram[1102]  = 0;
  ram[1103]  = 0;
  ram[1104]  = 0;
  ram[1105]  = 137;
  ram[1106]  = 255;
  ram[1107]  = 255;
  ram[1108]  = 255;
  ram[1109]  = 255;
  ram[1110]  = 255;
  ram[1111]  = 255;
  ram[1112]  = 255;
  ram[1113]  = 255;
  ram[1114]  = 255;
  ram[1115]  = 255;
  ram[1116]  = 255;
  ram[1117]  = 255;
  ram[1118]  = 255;
  ram[1119]  = 255;
  ram[1120]  = 255;
  ram[1121]  = 255;
  ram[1122]  = 255;
  ram[1123]  = 255;
  ram[1124]  = 255;
  ram[1125]  = 255;
  ram[1126]  = 255;
  ram[1127]  = 255;
  ram[1128]  = 255;
  ram[1129]  = 255;
  ram[1130]  = 255;
  ram[1131]  = 255;
  ram[1132]  = 137;
  ram[1133]  = 0;
  ram[1134]  = 0;
  ram[1135]  = 0;
  ram[1136]  = 0;
  ram[1137]  = 0;
  ram[1138]  = 0;
  ram[1139]  = 0;
  ram[1140]  = 0;
  ram[1141]  = 0;
  ram[1142]  = 0;
  ram[1143]  = 0;
  ram[1144]  = 0;
  ram[1145]  = 137;
  ram[1146]  = 255;
  ram[1147]  = 255;
  ram[1148]  = 255;
  ram[1149]  = 255;
  ram[1150]  = 255;
  ram[1151]  = 255;
  ram[1152]  = 255;
  ram[1153]  = 255;
  ram[1154]  = 255;
  ram[1155]  = 255;
  ram[1156]  = 255;
  ram[1157]  = 255;
  ram[1158]  = 255;
  ram[1159]  = 255;
  ram[1160]  = 255;
  ram[1161]  = 255;
  ram[1162]  = 255;
  ram[1163]  = 255;
  ram[1164]  = 255;
  ram[1165]  = 255;
  ram[1166]  = 255;
  ram[1167]  = 255;
  ram[1168]  = 255;
  ram[1169]  = 255;
  ram[1170]  = 255;
  ram[1171]  = 255;
  ram[1172]  = 255;
  ram[1173]  = 255;
  ram[1174]  = 255;
  ram[1175]  = 255;
  ram[1176]  = 255;
  ram[1177]  = 255;
  ram[1178]  = 255;
  ram[1179]  = 255;
  ram[1180]  = 255;
  ram[1181]  = 255;
  ram[1182]  = 255;
  ram[1183]  = 255;
  ram[1184]  = 255;
  ram[1185]  = 255;
  ram[1186]  = 255;
  ram[1187]  = 255;
  ram[1188]  = 255;
  ram[1189]  = 255;
  ram[1190]  = 255;
  ram[1191]  = 255;
  ram[1192]  = 255;
  ram[1193]  = 255;
  ram[1194]  = 255;
  ram[1195]  = 255;
  ram[1196]  = 255;
  ram[1197]  = 255;
  ram[1198]  = 255;
  ram[1199]  = 255;
  ram[1200]  = 255;
  ram[1201]  = 255;
  ram[1202]  = 255;
  ram[1203]  = 255;
  ram[1204]  = 255;
  ram[1205]  = 255;
  ram[1206]  = 255;
  ram[1207]  = 255;
  ram[1208]  = 255;
  ram[1209]  = 255;
  ram[1210]  = 255;
  ram[1211]  = 255;
  ram[1212]  = 255;
  ram[1213]  = 255;
  ram[1214]  = 255;
  ram[1215]  = 255;
  ram[1216]  = 255;
  ram[1217]  = 255;
  ram[1218]  = 255;
  ram[1219]  = 255;
  ram[1220]  = 255;
  ram[1221]  = 255;
  ram[1222]  = 255;
  ram[1223]  = 255;
  ram[1224]  = 255;
  ram[1225]  = 255;
  ram[1226]  = 255;
  ram[1227]  = 255;
  ram[1228]  = 255;
  ram[1229]  = 255;
  ram[1230]  = 255;
  ram[1231]  = 255;
  ram[1232]  = 255;
  ram[1233]  = 255;
  ram[1234]  = 255;
  ram[1235]  = 255;
  ram[1236]  = 255;
  ram[1237]  = 255;
  ram[1238]  = 255;
  ram[1239]  = 255;
  ram[1240]  = 255;
  ram[1241]  = 255;
  ram[1242]  = 255;
  ram[1243]  = 255;
  ram[1244]  = 255;
  ram[1245]  = 255;
  ram[1246]  = 255;
  ram[1247]  = 255;
  ram[1248]  = 255;
  ram[1249]  = 255;
  ram[1250]  = 255;
  ram[1251]  = 255;
  ram[1252]  = 255;
  ram[1253]  = 255;
  ram[1254]  = 255;
  ram[1255]  = 255;
  ram[1256]  = 255;
  ram[1257]  = 255;
  ram[1258]  = 255;
  ram[1259]  = 255;
  ram[1260]  = 255;
  ram[1261]  = 255;
  ram[1262]  = 255;
  ram[1263]  = 255;
  ram[1264]  = 255;
  ram[1265]  = 255;
  ram[1266]  = 255;
  ram[1267]  = 255;
  ram[1268]  = 255;
  ram[1269]  = 255;
  ram[1270]  = 255;
  ram[1271]  = 255;
  ram[1272]  = 255;
  ram[1273]  = 255;
  ram[1274]  = 255;
  ram[1275]  = 255;
  ram[1276]  = 255;
  ram[1277]  = 255;
  ram[1278]  = 255;
  ram[1279]  = 255;
  ram[1280]  = 255;
  ram[1281]  = 255;
  ram[1282]  = 255;
  ram[1283]  = 255;
  ram[1284]  = 255;
  ram[1285]  = 255;
  ram[1286]  = 255;
  ram[1287]  = 255;
  ram[1288]  = 255;
  ram[1289]  = 255;
  ram[1290]  = 255;
  ram[1291]  = 255;
  ram[1292]  = 255;
  ram[1293]  = 255;
  ram[1294]  = 255;
  ram[1295]  = 255;
  ram[1296]  = 255;
  ram[1297]  = 255;
  ram[1298]  = 255;
  ram[1299]  = 255;
  ram[1300]  = 255;
  ram[1301]  = 255;
  ram[1302]  = 255;
  ram[1303]  = 255;
  ram[1304]  = 255;
  ram[1305]  = 255;
  ram[1306]  = 255;
  ram[1307]  = 255;
  ram[1308]  = 255;
  ram[1309]  = 255;
  ram[1310]  = 255;
  ram[1311]  = 255;
  ram[1312]  = 255;
  ram[1313]  = 255;
  ram[1314]  = 255;
  ram[1315]  = 255;
  ram[1316]  = 255;
  ram[1317]  = 255;
  ram[1318]  = 255;
  ram[1319]  = 255;
  ram[1320]  = 255;
  ram[1321]  = 255;
  ram[1322]  = 255;
  ram[1323]  = 255;
  ram[1324]  = 255;
  ram[1325]  = 255;
  ram[1326]  = 255;
  ram[1327]  = 255;
  ram[1328]  = 255;
  ram[1329]  = 255;
  ram[1330]  = 255;
  ram[1331]  = 255;
  ram[1332]  = 255;
  ram[1333]  = 255;
  ram[1334]  = 255;
  ram[1335]  = 255;
  ram[1336]  = 255;
  ram[1337]  = 255;
  ram[1338]  = 255;
  ram[1339]  = 255;
  ram[1340]  = 255;
  ram[1341]  = 255;
  ram[1342]  = 255;
  ram[1343]  = 255;
  ram[1344]  = 255;
  ram[1345]  = 255;
  ram[1346]  = 255;
  ram[1347]  = 255;
  ram[1348]  = 255;
  ram[1349]  = 255;
  ram[1350]  = 255;
  ram[1351]  = 255;
  ram[1352]  = 255;
  ram[1353]  = 255;
  ram[1354]  = 255;
  ram[1355]  = 255;
  ram[1356]  = 255;
  ram[1357]  = 255;
  ram[1358]  = 255;
  ram[1359]  = 255;
  ram[1360]  = 255;
  ram[1361]  = 255;
  ram[1362]  = 255;
  ram[1363]  = 255;
  ram[1364]  = 255;
  ram[1365]  = 255;
  ram[1366]  = 255;
  ram[1367]  = 255;
  ram[1368]  = 255;
  ram[1369]  = 255;
  ram[1370]  = 255;
  ram[1371]  = 255;
  ram[1372]  = 255;
  ram[1373]  = 255;
  ram[1374]  = 255;
  ram[1375]  = 255;
  ram[1376]  = 255;
  ram[1377]  = 255;
  ram[1378]  = 255;
  ram[1379]  = 255;
  ram[1380]  = 255;
  ram[1381]  = 255;
  ram[1382]  = 255;
  ram[1383]  = 255;
  ram[1384]  = 255;
  ram[1385]  = 255;
  ram[1386]  = 255;
  ram[1387]  = 255;
  ram[1388]  = 255;
  ram[1389]  = 255;
  ram[1390]  = 255;
  ram[1391]  = 255;
  ram[1392]  = 255;
  ram[1393]  = 255;
  ram[1394]  = 255;
  ram[1395]  = 255;
  ram[1396]  = 255;
  ram[1397]  = 255;
  ram[1398]  = 255;
  ram[1399]  = 255;
  ram[1400]  = 255;
  ram[1401]  = 255;
  ram[1402]  = 255;
  ram[1403]  = 255;
  ram[1404]  = 255;
  ram[1405]  = 255;
  ram[1406]  = 255;
  ram[1407]  = 255;
  ram[1408]  = 255;
  ram[1409]  = 255;
  ram[1410]  = 255;
  ram[1411]  = 255;
  ram[1412]  = 255;
  ram[1413]  = 255;
  ram[1414]  = 255;
  ram[1415]  = 255;
  ram[1416]  = 255;
  ram[1417]  = 255;
  ram[1418]  = 255;
  ram[1419]  = 255;
  ram[1420]  = 255;
  ram[1421]  = 255;
  ram[1422]  = 255;
  ram[1423]  = 255;
  ram[1424]  = 255;
  ram[1425]  = 255;
  ram[1426]  = 255;
  ram[1427]  = 255;
  ram[1428]  = 255;
  ram[1429]  = 255;
  ram[1430]  = 255;
  ram[1431]  = 255;
  ram[1432]  = 255;
  ram[1433]  = 255;
  ram[1434]  = 255;
  ram[1435]  = 255;
  ram[1436]  = 255;
  ram[1437]  = 255;
  ram[1438]  = 255;
  ram[1439]  = 255;
  ram[1440]  = 255;
  ram[1441]  = 255;
  ram[1442]  = 255;
  ram[1443]  = 255;
  ram[1444]  = 255;
  ram[1445]  = 255;
  ram[1446]  = 255;
  ram[1447]  = 255;
  ram[1448]  = 255;
  ram[1449]  = 255;
  ram[1450]  = 255;
  ram[1451]  = 255;
  ram[1452]  = 255;
  ram[1453]  = 255;
  ram[1454]  = 255;
  ram[1455]  = 255;
  ram[1456]  = 255;
  ram[1457]  = 255;
  ram[1458]  = 255;
  ram[1459]  = 255;
  ram[1460]  = 255;
  ram[1461]  = 255;
  ram[1462]  = 255;
  ram[1463]  = 255;
  ram[1464]  = 255;
  ram[1465]  = 255;
  ram[1466]  = 255;
  ram[1467]  = 255;
  ram[1468]  = 255;
  ram[1469]  = 255;
  ram[1470]  = 255;
  ram[1471]  = 255;
  ram[1472]  = 255;
  ram[1473]  = 255;
  ram[1474]  = 255;
  ram[1475]  = 255;
  ram[1476]  = 255;
  ram[1477]  = 255;
  ram[1478]  = 255;
  ram[1479]  = 255;
  ram[1480]  = 255;
  ram[1481]  = 255;
  ram[1482]  = 255;
  ram[1483]  = 255;
  ram[1484]  = 255;
  ram[1485]  = 255;
  ram[1486]  = 255;
  ram[1487]  = 255;
  ram[1488]  = 255;
  ram[1489]  = 255;
  ram[1490]  = 255;
  ram[1491]  = 255;
  ram[1492]  = 255;
  ram[1493]  = 255;
  ram[1494]  = 255;
  ram[1495]  = 255;
  ram[1496]  = 255;
  ram[1497]  = 255;
  ram[1498]  = 255;
  ram[1499]  = 255;
  ram[1500]  = 255;
  ram[1501]  = 255;
  ram[1502]  = 255;
  ram[1503]  = 255;
  ram[1504]  = 255;
  ram[1505]  = 255;
  ram[1506]  = 255;
  ram[1507]  = 255;
  ram[1508]  = 255;
  ram[1509]  = 255;
  ram[1510]  = 255;
  ram[1511]  = 255;
  ram[1512]  = 255;
  ram[1513]  = 255;
  ram[1514]  = 255;
  ram[1515]  = 255;
  ram[1516]  = 255;
  ram[1517]  = 255;
  ram[1518]  = 255;
  ram[1519]  = 255;
  ram[1520]  = 255;
  ram[1521]  = 255;
  ram[1522]  = 255;
  ram[1523]  = 255;
  ram[1524]  = 255;
  ram[1525]  = 255;
  ram[1526]  = 255;
  ram[1527]  = 255;
  ram[1528]  = 255;
  ram[1529]  = 255;
  ram[1530]  = 255;
  ram[1531]  = 255;
  ram[1532]  = 255;
  ram[1533]  = 255;
  ram[1534]  = 255;
  ram[1535]  = 255;
  ram[1536]  = 255;
  ram[1537]  = 255;
  ram[1538]  = 255;
  ram[1539]  = 255;
  ram[1540]  = 255;
  ram[1541]  = 255;
  ram[1542]  = 255;
  ram[1543]  = 255;
  ram[1544]  = 255;
  ram[1545]  = 255;
  ram[1546]  = 255;
  ram[1547]  = 255;
  ram[1548]  = 255;
  ram[1549]  = 255;
  ram[1550]  = 255;
  ram[1551]  = 255;
  ram[1552]  = 255;
  ram[1553]  = 255;
  ram[1554]  = 255;
  ram[1555]  = 255;
  ram[1556]  = 255;
  ram[1557]  = 255;
  ram[1558]  = 255;
  ram[1559]  = 255;
  ram[1560]  = 255;
  ram[1561]  = 255;
  ram[1562]  = 255;
  ram[1563]  = 255;
  ram[1564]  = 255;
  ram[1565]  = 255;
  ram[1566]  = 255;
  ram[1567]  = 255;
  ram[1568]  = 255;
  ram[1569]  = 255;
  ram[1570]  = 255;
  ram[1571]  = 255;
  ram[1572]  = 255;
  ram[1573]  = 255;
  ram[1574]  = 255;
  ram[1575]  = 255;
  ram[1576]  = 255;
  ram[1577]  = 255;
  ram[1578]  = 255;
  ram[1579]  = 255;
  ram[1580]  = 255;
  ram[1581]  = 255;
  ram[1582]  = 255;
  ram[1583]  = 255;
  ram[1584]  = 255;
  ram[1585]  = 255;
  ram[1586]  = 255;
  ram[1587]  = 255;
  ram[1588]  = 255;
  ram[1589]  = 255;
  ram[1590]  = 255;
  ram[1591]  = 255;
  ram[1592]  = 255;
  ram[1593]  = 255;
  ram[1594]  = 255;
  ram[1595]  = 255;
  ram[1596]  = 255;
  ram[1597]  = 255;
  ram[1598]  = 255;
  ram[1599]  = 255;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
