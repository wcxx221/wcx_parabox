module rom_cai_r(clock, address, q);        // ROM-stored RGB bitmap for vegetable
input clock;
output [7:0] q;
input [8:0] address;
reg [7:0] dout;
reg [7:0] ram [511:0];
assign q = dout;

initial begin
  ram[0]  = 255;
  ram[1]  = 255;
  ram[2]  = 255;
  ram[3]  = 255;
  ram[4]  = 255;
  ram[5]  = 255;
  ram[6]  = 255;
  ram[7]  = 255;
  ram[8]  = 255;
  ram[9]  = 63;
  ram[10]  = 63;
  ram[11]  = 255;
  ram[12]  = 255;
  ram[13]  = 255;
  ram[14]  = 255;
  ram[15]  = 255;
  ram[16]  = 255;
  ram[17]  = 255;
  ram[18]  = 255;
  ram[19]  = 255;
  ram[20]  = 255;
  ram[21]  = 255;
  ram[22]  = 255;
  ram[23]  = 255;
  ram[24]  = 255;
  ram[25]  = 255;
  ram[26]  = 255;
  ram[27]  = 255;
  ram[28]  = 63;
  ram[29]  = 63;
  ram[30]  = 63;
  ram[31]  = 63;
  ram[32]  = 255;
  ram[33]  = 255;
  ram[34]  = 255;
  ram[35]  = 255;
  ram[36]  = 255;
  ram[37]  = 255;
  ram[38]  = 255;
  ram[39]  = 255;
  ram[40]  = 255;
  ram[41]  = 255;
  ram[42]  = 255;
  ram[43]  = 255;
  ram[44]  = 255;
  ram[45]  = 255;
  ram[46]  = 255;
  ram[47]  = 63;
  ram[48]  = 63;
  ram[49]  = 63;
  ram[50]  = 63;
  ram[51]  = 63;
  ram[52]  = 63;
  ram[53]  = 255;
  ram[54]  = 255;
  ram[55]  = 255;
  ram[56]  = 255;
  ram[57]  = 255;
  ram[58]  = 255;
  ram[59]  = 255;
  ram[60]  = 255;
  ram[61]  = 255;
  ram[62]  = 255;
  ram[63]  = 255;
  ram[64]  = 255;
  ram[65]  = 255;
  ram[66]  = 255;
  ram[67]  = 63;
  ram[68]  = 63;
  ram[69]  = 63;
  ram[70]  = 63;
  ram[71]  = 63;
  ram[72]  = 63;
  ram[73]  = 255;
  ram[74]  = 255;
  ram[75]  = 255;
  ram[76]  = 255;
  ram[77]  = 255;
  ram[78]  = 255;
  ram[79]  = 255;
  ram[80]  = 255;
  ram[81]  = 255;
  ram[82]  = 255;
  ram[83]  = 255;
  ram[84]  = 255;
  ram[85]  = 255;
  ram[86]  = 63;
  ram[87]  = 63;
  ram[88]  = 63;
  ram[89]  = 63;
  ram[90]  = 63;
  ram[91]  = 63;
  ram[92]  = 63;
  ram[93]  = 63;
  ram[94]  = 255;
  ram[95]  = 255;
  ram[96]  = 255;
  ram[97]  = 255;
  ram[98]  = 255;
  ram[99]  = 255;
  ram[100]  = 255;
  ram[101]  = 255;
  ram[102]  = 255;
  ram[103]  = 255;
  ram[104]  = 255;
  ram[105]  = 255;
  ram[106]  = 63;
  ram[107]  = 63;
  ram[108]  = 63;
  ram[109]  = 63;
  ram[110]  = 63;
  ram[111]  = 63;
  ram[112]  = 63;
  ram[113]  = 63;
  ram[114]  = 255;
  ram[115]  = 255;
  ram[116]  = 255;
  ram[117]  = 255;
  ram[118]  = 255;
  ram[119]  = 255;
  ram[120]  = 255;
  ram[121]  = 255;
  ram[122]  = 255;
  ram[123]  = 255;
  ram[124]  = 255;
  ram[125]  = 63;
  ram[126]  = 63;
  ram[127]  = 63;
  ram[128]  = 63;
  ram[129]  = 63;
  ram[130]  = 63;
  ram[131]  = 63;
  ram[132]  = 63;
  ram[133]  = 63;
  ram[134]  = 63;
  ram[135]  = 255;
  ram[136]  = 255;
  ram[137]  = 255;
  ram[138]  = 255;
  ram[139]  = 255;
  ram[140]  = 255;
  ram[141]  = 255;
  ram[142]  = 255;
  ram[143]  = 255;
  ram[144]  = 255;
  ram[145]  = 63;
  ram[146]  = 63;
  ram[147]  = 63;
  ram[148]  = 63;
  ram[149]  = 63;
  ram[150]  = 63;
  ram[151]  = 63;
  ram[152]  = 63;
  ram[153]  = 63;
  ram[154]  = 63;
  ram[155]  = 255;
  ram[156]  = 255;
  ram[157]  = 255;
  ram[158]  = 255;
  ram[159]  = 255;
  ram[160]  = 255;
  ram[161]  = 255;
  ram[162]  = 255;
  ram[163]  = 255;
  ram[164]  = 63;
  ram[165]  = 63;
  ram[166]  = 63;
  ram[167]  = 63;
  ram[168]  = 63;
  ram[169]  = 63;
  ram[170]  = 63;
  ram[171]  = 63;
  ram[172]  = 63;
  ram[173]  = 63;
  ram[174]  = 63;
  ram[175]  = 63;
  ram[176]  = 255;
  ram[177]  = 255;
  ram[178]  = 255;
  ram[179]  = 255;
  ram[180]  = 255;
  ram[181]  = 255;
  ram[182]  = 255;
  ram[183]  = 255;
  ram[184]  = 63;
  ram[185]  = 63;
  ram[186]  = 63;
  ram[187]  = 63;
  ram[188]  = 63;
  ram[189]  = 255;
  ram[190]  = 255;
  ram[191]  = 63;
  ram[192]  = 63;
  ram[193]  = 63;
  ram[194]  = 63;
  ram[195]  = 63;
  ram[196]  = 255;
  ram[197]  = 255;
  ram[198]  = 255;
  ram[199]  = 255;
  ram[200]  = 255;
  ram[201]  = 255;
  ram[202]  = 255;
  ram[203]  = 63;
  ram[204]  = 63;
  ram[205]  = 63;
  ram[206]  = 63;
  ram[207]  = 63;
  ram[208]  = 63;
  ram[209]  = 255;
  ram[210]  = 255;
  ram[211]  = 63;
  ram[212]  = 63;
  ram[213]  = 63;
  ram[214]  = 63;
  ram[215]  = 63;
  ram[216]  = 63;
  ram[217]  = 255;
  ram[218]  = 255;
  ram[219]  = 255;
  ram[220]  = 255;
  ram[221]  = 255;
  ram[222]  = 255;
  ram[223]  = 63;
  ram[224]  = 63;
  ram[225]  = 63;
  ram[226]  = 63;
  ram[227]  = 63;
  ram[228]  = 255;
  ram[229]  = 255;
  ram[230]  = 255;
  ram[231]  = 255;
  ram[232]  = 63;
  ram[233]  = 63;
  ram[234]  = 63;
  ram[235]  = 63;
  ram[236]  = 63;
  ram[237]  = 255;
  ram[238]  = 255;
  ram[239]  = 255;
  ram[240]  = 255;
  ram[241]  = 255;
  ram[242]  = 63;
  ram[243]  = 63;
  ram[244]  = 63;
  ram[245]  = 63;
  ram[246]  = 63;
  ram[247]  = 63;
  ram[248]  = 255;
  ram[249]  = 255;
  ram[250]  = 255;
  ram[251]  = 255;
  ram[252]  = 63;
  ram[253]  = 63;
  ram[254]  = 63;
  ram[255]  = 63;
  ram[256]  = 63;
  ram[257]  = 63;
  ram[258]  = 255;
  ram[259]  = 255;
  ram[260]  = 255;
  ram[261]  = 255;
  ram[262]  = 63;
  ram[263]  = 63;
  ram[264]  = 63;
  ram[265]  = 63;
  ram[266]  = 63;
  ram[267]  = 255;
  ram[268]  = 255;
  ram[269]  = 255;
  ram[270]  = 255;
  ram[271]  = 255;
  ram[272]  = 255;
  ram[273]  = 63;
  ram[274]  = 63;
  ram[275]  = 63;
  ram[276]  = 63;
  ram[277]  = 63;
  ram[278]  = 255;
  ram[279]  = 255;
  ram[280]  = 255;
  ram[281]  = 63;
  ram[282]  = 63;
  ram[283]  = 63;
  ram[284]  = 63;
  ram[285]  = 63;
  ram[286]  = 63;
  ram[287]  = 255;
  ram[288]  = 255;
  ram[289]  = 255;
  ram[290]  = 255;
  ram[291]  = 255;
  ram[292]  = 255;
  ram[293]  = 63;
  ram[294]  = 63;
  ram[295]  = 63;
  ram[296]  = 63;
  ram[297]  = 63;
  ram[298]  = 63;
  ram[299]  = 255;
  ram[300]  = 255;
  ram[301]  = 63;
  ram[302]  = 63;
  ram[303]  = 63;
  ram[304]  = 63;
  ram[305]  = 63;
  ram[306]  = 63;
  ram[307]  = 63;
  ram[308]  = 63;
  ram[309]  = 63;
  ram[310]  = 63;
  ram[311]  = 63;
  ram[312]  = 63;
  ram[313]  = 63;
  ram[314]  = 63;
  ram[315]  = 63;
  ram[316]  = 63;
  ram[317]  = 63;
  ram[318]  = 63;
  ram[319]  = 255;
  ram[320]  = 63;
  ram[321]  = 63;
  ram[322]  = 63;
  ram[323]  = 63;
  ram[324]  = 63;
  ram[325]  = 63;
  ram[326]  = 63;
  ram[327]  = 63;
  ram[328]  = 63;
  ram[329]  = 63;
  ram[330]  = 63;
  ram[331]  = 63;
  ram[332]  = 63;
  ram[333]  = 63;
  ram[334]  = 63;
  ram[335]  = 63;
  ram[336]  = 63;
  ram[337]  = 63;
  ram[338]  = 63;
  ram[339]  = 63;
  ram[340]  = 63;
  ram[341]  = 63;
  ram[342]  = 63;
  ram[343]  = 63;
  ram[344]  = 63;
  ram[345]  = 63;
  ram[346]  = 63;
  ram[347]  = 63;
  ram[348]  = 63;
  ram[349]  = 63;
  ram[350]  = 63;
  ram[351]  = 63;
  ram[352]  = 63;
  ram[353]  = 63;
  ram[354]  = 63;
  ram[355]  = 63;
  ram[356]  = 63;
  ram[357]  = 63;
  ram[358]  = 63;
  ram[359]  = 63;
  ram[360]  = 63;
  ram[361]  = 63;
  ram[362]  = 63;
  ram[363]  = 63;
  ram[364]  = 63;
  ram[365]  = 63;
  ram[366]  = 63;
  ram[367]  = 63;
  ram[368]  = 63;
  ram[369]  = 63;
  ram[370]  = 63;
  ram[371]  = 63;
  ram[372]  = 63;
  ram[373]  = 63;
  ram[374]  = 63;
  ram[375]  = 63;
  ram[376]  = 63;
  ram[377]  = 63;
  ram[378]  = 63;
  ram[379]  = 63;
  ram[380]  = 255;
  ram[381]  = 63;
  ram[382]  = 63;
  ram[383]  = 63;
  ram[384]  = 63;
  ram[385]  = 63;
  ram[386]  = 63;
  ram[387]  = 63;
  ram[388]  = 63;
  ram[389]  = 63;
  ram[390]  = 63;
  ram[391]  = 63;
  ram[392]  = 63;
  ram[393]  = 63;
  ram[394]  = 63;
  ram[395]  = 63;
  ram[396]  = 63;
  ram[397]  = 63;
  ram[398]  = 63;
  ram[399]  = 255;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
