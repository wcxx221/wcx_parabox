module rom_cai_b(clock, address, q);        // ROM-stored RGB bitmap for cai
input clock;
output [7:0] q;
input [8:0] address;
reg [7:0] dout;
reg [7:0] ram [511:0];
assign q = dout;

initial begin
  ram[0]  = 255;
  ram[1]  = 255;
  ram[2]  = 255;
  ram[3]  = 255;
  ram[4]  = 255;
  ram[5]  = 255;
  ram[6]  = 255;
  ram[7]  = 255;
  ram[8]  = 255;
  ram[9]  = 204;
  ram[10]  = 204;
  ram[11]  = 255;
  ram[12]  = 255;
  ram[13]  = 255;
  ram[14]  = 255;
  ram[15]  = 255;
  ram[16]  = 255;
  ram[17]  = 255;
  ram[18]  = 255;
  ram[19]  = 255;
  ram[20]  = 255;
  ram[21]  = 255;
  ram[22]  = 255;
  ram[23]  = 255;
  ram[24]  = 255;
  ram[25]  = 255;
  ram[26]  = 255;
  ram[27]  = 255;
  ram[28]  = 204;
  ram[29]  = 204;
  ram[30]  = 204;
  ram[31]  = 204;
  ram[32]  = 255;
  ram[33]  = 255;
  ram[34]  = 255;
  ram[35]  = 255;
  ram[36]  = 255;
  ram[37]  = 255;
  ram[38]  = 255;
  ram[39]  = 255;
  ram[40]  = 255;
  ram[41]  = 255;
  ram[42]  = 255;
  ram[43]  = 255;
  ram[44]  = 255;
  ram[45]  = 255;
  ram[46]  = 255;
  ram[47]  = 204;
  ram[48]  = 204;
  ram[49]  = 204;
  ram[50]  = 204;
  ram[51]  = 204;
  ram[52]  = 204;
  ram[53]  = 255;
  ram[54]  = 255;
  ram[55]  = 255;
  ram[56]  = 255;
  ram[57]  = 255;
  ram[58]  = 255;
  ram[59]  = 255;
  ram[60]  = 255;
  ram[61]  = 255;
  ram[62]  = 255;
  ram[63]  = 255;
  ram[64]  = 255;
  ram[65]  = 255;
  ram[66]  = 255;
  ram[67]  = 204;
  ram[68]  = 204;
  ram[69]  = 204;
  ram[70]  = 204;
  ram[71]  = 204;
  ram[72]  = 204;
  ram[73]  = 255;
  ram[74]  = 255;
  ram[75]  = 255;
  ram[76]  = 255;
  ram[77]  = 255;
  ram[78]  = 255;
  ram[79]  = 255;
  ram[80]  = 255;
  ram[81]  = 255;
  ram[82]  = 255;
  ram[83]  = 255;
  ram[84]  = 255;
  ram[85]  = 255;
  ram[86]  = 204;
  ram[87]  = 204;
  ram[88]  = 204;
  ram[89]  = 204;
  ram[90]  = 204;
  ram[91]  = 204;
  ram[92]  = 204;
  ram[93]  = 204;
  ram[94]  = 255;
  ram[95]  = 255;
  ram[96]  = 255;
  ram[97]  = 255;
  ram[98]  = 255;
  ram[99]  = 255;
  ram[100]  = 255;
  ram[101]  = 255;
  ram[102]  = 255;
  ram[103]  = 255;
  ram[104]  = 255;
  ram[105]  = 255;
  ram[106]  = 204;
  ram[107]  = 204;
  ram[108]  = 204;
  ram[109]  = 204;
  ram[110]  = 204;
  ram[111]  = 204;
  ram[112]  = 204;
  ram[113]  = 204;
  ram[114]  = 255;
  ram[115]  = 255;
  ram[116]  = 255;
  ram[117]  = 255;
  ram[118]  = 255;
  ram[119]  = 255;
  ram[120]  = 255;
  ram[121]  = 255;
  ram[122]  = 255;
  ram[123]  = 255;
  ram[124]  = 255;
  ram[125]  = 204;
  ram[126]  = 204;
  ram[127]  = 204;
  ram[128]  = 204;
  ram[129]  = 204;
  ram[130]  = 204;
  ram[131]  = 204;
  ram[132]  = 204;
  ram[133]  = 204;
  ram[134]  = 204;
  ram[135]  = 255;
  ram[136]  = 255;
  ram[137]  = 255;
  ram[138]  = 255;
  ram[139]  = 255;
  ram[140]  = 255;
  ram[141]  = 255;
  ram[142]  = 255;
  ram[143]  = 255;
  ram[144]  = 255;
  ram[145]  = 204;
  ram[146]  = 204;
  ram[147]  = 204;
  ram[148]  = 204;
  ram[149]  = 204;
  ram[150]  = 204;
  ram[151]  = 204;
  ram[152]  = 204;
  ram[153]  = 204;
  ram[154]  = 204;
  ram[155]  = 255;
  ram[156]  = 255;
  ram[157]  = 255;
  ram[158]  = 255;
  ram[159]  = 255;
  ram[160]  = 255;
  ram[161]  = 255;
  ram[162]  = 255;
  ram[163]  = 255;
  ram[164]  = 204;
  ram[165]  = 204;
  ram[166]  = 204;
  ram[167]  = 204;
  ram[168]  = 204;
  ram[169]  = 204;
  ram[170]  = 204;
  ram[171]  = 204;
  ram[172]  = 204;
  ram[173]  = 204;
  ram[174]  = 204;
  ram[175]  = 204;
  ram[176]  = 255;
  ram[177]  = 255;
  ram[178]  = 255;
  ram[179]  = 255;
  ram[180]  = 255;
  ram[181]  = 255;
  ram[182]  = 255;
  ram[183]  = 255;
  ram[184]  = 204;
  ram[185]  = 204;
  ram[186]  = 204;
  ram[187]  = 204;
  ram[188]  = 204;
  ram[189]  = 255;
  ram[190]  = 255;
  ram[191]  = 204;
  ram[192]  = 204;
  ram[193]  = 204;
  ram[194]  = 204;
  ram[195]  = 204;
  ram[196]  = 255;
  ram[197]  = 255;
  ram[198]  = 255;
  ram[199]  = 255;
  ram[200]  = 255;
  ram[201]  = 255;
  ram[202]  = 255;
  ram[203]  = 204;
  ram[204]  = 204;
  ram[205]  = 204;
  ram[206]  = 204;
  ram[207]  = 204;
  ram[208]  = 204;
  ram[209]  = 255;
  ram[210]  = 255;
  ram[211]  = 204;
  ram[212]  = 204;
  ram[213]  = 204;
  ram[214]  = 204;
  ram[215]  = 204;
  ram[216]  = 204;
  ram[217]  = 255;
  ram[218]  = 255;
  ram[219]  = 255;
  ram[220]  = 255;
  ram[221]  = 255;
  ram[222]  = 255;
  ram[223]  = 204;
  ram[224]  = 204;
  ram[225]  = 204;
  ram[226]  = 204;
  ram[227]  = 204;
  ram[228]  = 255;
  ram[229]  = 255;
  ram[230]  = 255;
  ram[231]  = 255;
  ram[232]  = 204;
  ram[233]  = 204;
  ram[234]  = 204;
  ram[235]  = 204;
  ram[236]  = 204;
  ram[237]  = 255;
  ram[238]  = 255;
  ram[239]  = 255;
  ram[240]  = 255;
  ram[241]  = 255;
  ram[242]  = 204;
  ram[243]  = 204;
  ram[244]  = 204;
  ram[245]  = 204;
  ram[246]  = 204;
  ram[247]  = 204;
  ram[248]  = 255;
  ram[249]  = 255;
  ram[250]  = 255;
  ram[251]  = 255;
  ram[252]  = 204;
  ram[253]  = 204;
  ram[254]  = 204;
  ram[255]  = 204;
  ram[256]  = 204;
  ram[257]  = 204;
  ram[258]  = 255;
  ram[259]  = 255;
  ram[260]  = 255;
  ram[261]  = 255;
  ram[262]  = 204;
  ram[263]  = 204;
  ram[264]  = 204;
  ram[265]  = 204;
  ram[266]  = 204;
  ram[267]  = 255;
  ram[268]  = 255;
  ram[269]  = 255;
  ram[270]  = 255;
  ram[271]  = 255;
  ram[272]  = 255;
  ram[273]  = 204;
  ram[274]  = 204;
  ram[275]  = 204;
  ram[276]  = 204;
  ram[277]  = 204;
  ram[278]  = 255;
  ram[279]  = 255;
  ram[280]  = 255;
  ram[281]  = 204;
  ram[282]  = 204;
  ram[283]  = 204;
  ram[284]  = 204;
  ram[285]  = 204;
  ram[286]  = 204;
  ram[287]  = 255;
  ram[288]  = 255;
  ram[289]  = 255;
  ram[290]  = 255;
  ram[291]  = 255;
  ram[292]  = 255;
  ram[293]  = 204;
  ram[294]  = 204;
  ram[295]  = 204;
  ram[296]  = 204;
  ram[297]  = 204;
  ram[298]  = 204;
  ram[299]  = 255;
  ram[300]  = 255;
  ram[301]  = 204;
  ram[302]  = 204;
  ram[303]  = 204;
  ram[304]  = 204;
  ram[305]  = 204;
  ram[306]  = 204;
  ram[307]  = 204;
  ram[308]  = 204;
  ram[309]  = 204;
  ram[310]  = 204;
  ram[311]  = 204;
  ram[312]  = 204;
  ram[313]  = 204;
  ram[314]  = 204;
  ram[315]  = 204;
  ram[316]  = 204;
  ram[317]  = 204;
  ram[318]  = 204;
  ram[319]  = 255;
  ram[320]  = 204;
  ram[321]  = 204;
  ram[322]  = 204;
  ram[323]  = 204;
  ram[324]  = 204;
  ram[325]  = 204;
  ram[326]  = 204;
  ram[327]  = 204;
  ram[328]  = 204;
  ram[329]  = 204;
  ram[330]  = 204;
  ram[331]  = 204;
  ram[332]  = 204;
  ram[333]  = 204;
  ram[334]  = 204;
  ram[335]  = 204;
  ram[336]  = 204;
  ram[337]  = 204;
  ram[338]  = 204;
  ram[339]  = 204;
  ram[340]  = 204;
  ram[341]  = 204;
  ram[342]  = 204;
  ram[343]  = 204;
  ram[344]  = 204;
  ram[345]  = 204;
  ram[346]  = 204;
  ram[347]  = 204;
  ram[348]  = 204;
  ram[349]  = 204;
  ram[350]  = 204;
  ram[351]  = 204;
  ram[352]  = 204;
  ram[353]  = 204;
  ram[354]  = 204;
  ram[355]  = 204;
  ram[356]  = 204;
  ram[357]  = 204;
  ram[358]  = 204;
  ram[359]  = 204;
  ram[360]  = 204;
  ram[361]  = 204;
  ram[362]  = 204;
  ram[363]  = 204;
  ram[364]  = 204;
  ram[365]  = 204;
  ram[366]  = 204;
  ram[367]  = 204;
  ram[368]  = 204;
  ram[369]  = 204;
  ram[370]  = 204;
  ram[371]  = 204;
  ram[372]  = 204;
  ram[373]  = 204;
  ram[374]  = 204;
  ram[375]  = 204;
  ram[376]  = 204;
  ram[377]  = 204;
  ram[378]  = 204;
  ram[379]  = 204;
  ram[380]  = 255;
  ram[381]  = 204;
  ram[382]  = 204;
  ram[383]  = 204;
  ram[384]  = 204;
  ram[385]  = 204;
  ram[386]  = 204;
  ram[387]  = 204;
  ram[388]  = 204;
  ram[389]  = 204;
  ram[390]  = 204;
  ram[391]  = 204;
  ram[392]  = 204;
  ram[393]  = 204;
  ram[394]  = 204;
  ram[395]  = 204;
  ram[396]  = 204;
  ram[397]  = 204;
  ram[398]  = 204;
  ram[399]  = 255;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
