module rom_man_b(clock, address, q);        // ROM-stored RGB bitmap for player(man)
input clock;
output [7:0] q;
input [8:0] address;
reg [7:0] dout;
reg [7:0] ram [511:0];
assign q = dout;

initial begin
  ram[0]  = 149;
  ram[1]  = 147;
  ram[2]  = 141;
  ram[3]  = 145;
  ram[4]  = 151;
  ram[5]  = 149;
  ram[6]  = 146;
  ram[7]  = 145;
  ram[8]  = 135;
  ram[9]  = 123;
  ram[10]  = 133;
  ram[11]  = 143;
  ram[12]  = 146;
  ram[13]  = 151;
  ram[14]  = 149;
  ram[15]  = 147;
  ram[16]  = 149;
  ram[17]  = 146;
  ram[18]  = 142;
  ram[19]  = 204;
  ram[20]  = 145;
  ram[21]  = 146;
  ram[22]  = 149;
  ram[23]  = 152;
  ram[24]  = 131;
  ram[25]  = 101;
  ram[26]  = 82;
  ram[27]  = 69;
  ram[28]  = 70;
  ram[29]  = 74;
  ram[30]  = 74;
  ram[31]  = 67;
  ram[32]  = 82;
  ram[33]  = 92;
  ram[34]  = 110;
  ram[35]  = 135;
  ram[36]  = 147;
  ram[37]  = 145;
  ram[38]  = 143;
  ram[39]  = 179;
  ram[40]  = 146;
  ram[41]  = 143;
  ram[42]  = 142;
  ram[43]  = 114;
  ram[44]  = 66;
  ram[45]  = 40;
  ram[46]  = 38;
  ram[47]  = 38;
  ram[48]  = 54;
  ram[49]  = 65;
  ram[50]  = 57;
  ram[51]  = 41;
  ram[52]  = 38;
  ram[53]  = 39;
  ram[54]  = 53;
  ram[55]  = 97;
  ram[56]  = 145;
  ram[57]  = 152;
  ram[58]  = 144;
  ram[59]  = 177;
  ram[60]  = 152;
  ram[61]  = 145;
  ram[62]  = 104;
  ram[63]  = 58;
  ram[64]  = 40;
  ram[65]  = 39;
  ram[66]  = 40;
  ram[67]  = 42;
  ram[68]  = 58;
  ram[69]  = 66;
  ram[70]  = 64;
  ram[71]  = 47;
  ram[72]  = 40;
  ram[73]  = 40;
  ram[74]  = 38;
  ram[75]  = 49;
  ram[76]  = 93;
  ram[77]  = 137;
  ram[78]  = 146;
  ram[79]  = 178;
  ram[80]  = 151;
  ram[81]  = 125;
  ram[82]  = 67;
  ram[83]  = 39;
  ram[84]  = 40;
  ram[85]  = 42;
  ram[86]  = 40;
  ram[87]  = 46;
  ram[88]  = 63;
  ram[89]  = 65;
  ram[90]  = 64;
  ram[91]  = 52;
  ram[92]  = 41;
  ram[93]  = 41;
  ram[94]  = 41;
  ram[95]  = 38;
  ram[96]  = 51;
  ram[97]  = 101;
  ram[98]  = 142;
  ram[99]  = 178;
  ram[100]  = 145;
  ram[101]  = 94;
  ram[102]  = 49;
  ram[103]  = 39;
  ram[104]  = 42;
  ram[105]  = 42;
  ram[106]  = 41;
  ram[107]  = 50;
  ram[108]  = 64;
  ram[109]  = 64;
  ram[110]  = 62;
  ram[111]  = 55;
  ram[112]  = 44;
  ram[113]  = 41;
  ram[114]  = 41;
  ram[115]  = 41;
  ram[116]  = 42;
  ram[117]  = 70;
  ram[118]  = 123;
  ram[119]  = 180;
  ram[120]  = 139;
  ram[121]  = 80;
  ram[122]  = 44;
  ram[123]  = 41;
  ram[124]  = 41;
  ram[125]  = 40;
  ram[126]  = 42;
  ram[127]  = 56;
  ram[128]  = 62;
  ram[129]  = 56;
  ram[130]  = 54;
  ram[131]  = 59;
  ram[132]  = 45;
  ram[133]  = 39;
  ram[134]  = 40;
  ram[135]  = 42;
  ram[136]  = 41;
  ram[137]  = 50;
  ram[138]  = 110;
  ram[139]  = 180;
  ram[140]  = 136;
  ram[141]  = 82;
  ram[142]  = 42;
  ram[143]  = 36;
  ram[144]  = 30;
  ram[145]  = 33;
  ram[146]  = 36;
  ram[147]  = 42;
  ram[148]  = 58;
  ram[149]  = 60;
  ram[150]  = 51;
  ram[151]  = 42;
  ram[152]  = 38;
  ram[153]  = 37;
  ram[154]  = 30;
  ram[155]  = 33;
  ram[156]  = 36;
  ram[157]  = 52;
  ram[158]  = 110;
  ram[159]  = 179;
  ram[160]  = 139;
  ram[161]  = 81;
  ram[162]  = 34;
  ram[163]  = 32;
  ram[164]  = 77;
  ram[165]  = 113;
  ram[166]  = 51;
  ram[167]  = 39;
  ram[168]  = 135;
  ram[169]  = 197;
  ram[170]  = 151;
  ram[171]  = 53;
  ram[172]  = 45;
  ram[173]  = 115;
  ram[174]  = 127;
  ram[175]  = 60;
  ram[176]  = 28;
  ram[177]  = 45;
  ram[178]  = 104;
  ram[179]  = 177;
  ram[180]  = 139;
  ram[181]  = 89;
  ram[182]  = 34;
  ram[183]  = 88;
  ram[184]  = 193;
  ram[185]  = 166;
  ram[186]  = 58;
  ram[187]  = 45;
  ram[188]  = 127;
  ram[189]  = 217;
  ram[190]  = 164;
  ram[191]  = 58;
  ram[192]  = 47;
  ram[193]  = 134;
  ram[194]  = 215;
  ram[195]  = 168;
  ram[196]  = 59;
  ram[197]  = 51;
  ram[198]  = 114;
  ram[199]  = 178;
  ram[200]  = 148;
  ram[201]  = 140;
  ram[202]  = 108;
  ram[203]  = 132;
  ram[204]  = 207;
  ram[205]  = 185;
  ram[206]  = 70;
  ram[207]  = 41;
  ram[208]  = 150;
  ram[209]  = 206;
  ram[210]  = 178;
  ram[211]  = 67;
  ram[212]  = 50;
  ram[213]  = 160;
  ram[214]  = 214;
  ram[215]  = 185;
  ram[216]  = 113;
  ram[217]  = 121;
  ram[218]  = 138;
  ram[219]  = 176;
  ram[220]  = 138;
  ram[221]  = 149;
  ram[222]  = 153;
  ram[223]  = 136;
  ram[224]  = 170;
  ram[225]  = 206;
  ram[226]  = 160;
  ram[227]  = 143;
  ram[228]  = 195;
  ram[229]  = 198;
  ram[230]  = 199;
  ram[231]  = 161;
  ram[232]  = 149;
  ram[233]  = 200;
  ram[234]  = 196;
  ram[235]  = 154;
  ram[236]  = 143;
  ram[237]  = 151;
  ram[238]  = 148;
  ram[239]  = 178;
  ram[240]  = 141;
  ram[241]  = 142;
  ram[242]  = 149;
  ram[243]  = 163;
  ram[244]  = 169;
  ram[245]  = 188;
  ram[246]  = 196;
  ram[247]  = 201;
  ram[248]  = 196;
  ram[249]  = 189;
  ram[250]  = 191;
  ram[251]  = 197;
  ram[252]  = 198;
  ram[253]  = 194;
  ram[254]  = 169;
  ram[255]  = 167;
  ram[256]  = 155;
  ram[257]  = 142;
  ram[258]  = 145;
  ram[259]  = 178;
  ram[260]  = 150;
  ram[261]  = 151;
  ram[262]  = 160;
  ram[263]  = 169;
  ram[264]  = 173;
  ram[265]  = 176;
  ram[266]  = 190;
  ram[267]  = 200;
  ram[268]  = 191;
  ram[269]  = 188;
  ram[270]  = 190;
  ram[271]  = 195;
  ram[272]  = 199;
  ram[273]  = 185;
  ram[274]  = 165;
  ram[275]  = 168;
  ram[276]  = 170;
  ram[277]  = 149;
  ram[278]  = 143;
  ram[279]  = 177;
  ram[280]  = 147;
  ram[281]  = 150;
  ram[282]  = 160;
  ram[283]  = 167;
  ram[284]  = 165;
  ram[285]  = 177;
  ram[286]  = 185;
  ram[287]  = 188;
  ram[288]  = 188;
  ram[289]  = 188;
  ram[290]  = 192;
  ram[291]  = 189;
  ram[292]  = 186;
  ram[293]  = 183;
  ram[294]  = 165;
  ram[295]  = 165;
  ram[296]  = 169;
  ram[297]  = 151;
  ram[298]  = 143;
  ram[299]  = 177;
  ram[300]  = 143;
  ram[301]  = 140;
  ram[302]  = 155;
  ram[303]  = 194;
  ram[304]  = 192;
  ram[305]  = 181;
  ram[306]  = 187;
  ram[307]  = 192;
  ram[308]  = 189;
  ram[309]  = 188;
  ram[310]  = 191;
  ram[311]  = 191;
  ram[312]  = 191;
  ram[313]  = 182;
  ram[314]  = 176;
  ram[315]  = 202;
  ram[316]  = 187;
  ram[317]  = 143;
  ram[318]  = 143;
  ram[319]  = 178;
  ram[320]  = 142;
  ram[321]  = 144;
  ram[322]  = 154;
  ram[323]  = 206;
  ram[324]  = 208;
  ram[325]  = 187;
  ram[326]  = 184;
  ram[327]  = 187;
  ram[328]  = 191;
  ram[329]  = 194;
  ram[330]  = 192;
  ram[331]  = 191;
  ram[332]  = 189;
  ram[333]  = 186;
  ram[334]  = 196;
  ram[335]  = 210;
  ram[336]  = 181;
  ram[337]  = 136;
  ram[338]  = 142;
  ram[339]  = 178;
  ram[340]  = 147;
  ram[341]  = 151;
  ram[342]  = 143;
  ram[343]  = 152;
  ram[344]  = 152;
  ram[345]  = 139;
  ram[346]  = 124;
  ram[347]  = 106;
  ram[348]  = 124;
  ram[349]  = 182;
  ram[350]  = 162;
  ram[351]  = 109;
  ram[352]  = 111;
  ram[353]  = 134;
  ram[354]  = 148;
  ram[355]  = 155;
  ram[356]  = 147;
  ram[357]  = 145;
  ram[358]  = 143;
  ram[359]  = 177;
  ram[360]  = 147;
  ram[361]  = 151;
  ram[362]  = 147;
  ram[363]  = 141;
  ram[364]  = 138;
  ram[365]  = 118;
  ram[366]  = 72;
  ram[367]  = 59;
  ram[368]  = 70;
  ram[369]  = 123;
  ram[370]  = 104;
  ram[371]  = 65;
  ram[372]  = 68;
  ram[373]  = 88;
  ram[374]  = 131;
  ram[375]  = 146;
  ram[376]  = 149;
  ram[377]  = 147;
  ram[378]  = 144;
  ram[379]  = 178;
  ram[380]  = 146;
  ram[381]  = 149;
  ram[382]  = 147;
  ram[383]  = 145;
  ram[384]  = 146;
  ram[385]  = 143;
  ram[386]  = 128;
  ram[387]  = 120;
  ram[388]  = 118;
  ram[389]  = 134;
  ram[390]  = 131;
  ram[391]  = 123;
  ram[392]  = 122;
  ram[393]  = 128;
  ram[394]  = 141;
  ram[395]  = 146;
  ram[396]  = 146;
  ram[397]  = 144;
  ram[398]  = 144;
  ram[399]  = 178;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
