module rom_dist_r(clock, address, q);  // ROM-stored RGB bitmap for level destination
input clock;
output [7:0] q;
input [8:0] address;
reg [7:0] dout;
reg [7:0] ram [511:0];
assign q = dout;
        //Simple synchronous ROM module storing 8-bit pixel data
initial begin
  ram[0]  = 255;
  ram[1]  = 255;
  ram[2]  = 255;
  ram[3]  = 255;
  ram[4]  = 255;
  ram[5]  = 255;
  ram[6]  = 255;
  ram[7]  = 232;
  ram[8]  = 232;
  ram[9]  = 232;
  ram[10]  = 232;
  ram[11]  = 232;
  ram[12]  = 255;
  ram[13]  = 255;
  ram[14]  = 255;
  ram[15]  = 255;
  ram[16]  = 255;
  ram[17]  = 255;
  ram[18]  = 255;
  ram[19]  = 255;
  ram[20]  = 255;
  ram[21]  = 255;
  ram[22]  = 255;
  ram[23]  = 255;
  ram[24]  = 255;
  ram[25]  = 232;
  ram[26]  = 232;
  ram[27]  = 232;
  ram[28]  = 232;
  ram[29]  = 232;
  ram[30]  = 232;
  ram[31]  = 232;
  ram[32]  = 232;
  ram[33]  = 232;
  ram[34]  = 255;
  ram[35]  = 255;
  ram[36]  = 255;
  ram[37]  = 255;
  ram[38]  = 255;
  ram[39]  = 255;
  ram[40]  = 255;
  ram[41]  = 255;
  ram[42]  = 255;
  ram[43]  = 232;
  ram[44]  = 232;
  ram[45]  = 232;
  ram[46]  = 232;
  ram[47]  = 232;
  ram[48]  = 232;
  ram[49]  = 232;
  ram[50]  = 232;
  ram[51]  = 232;
  ram[52]  = 232;
  ram[53]  = 232;
  ram[54]  = 232;
  ram[55]  = 232;
  ram[56]  = 255;
  ram[57]  = 255;
  ram[58]  = 255;
  ram[59]  = 255;
  ram[60]  = 255;
  ram[61]  = 255;
  ram[62]  = 232;
  ram[63]  = 232;
  ram[64]  = 232;
  ram[65]  = 232;
  ram[66]  = 232;
  ram[67]  = 232;
  ram[68]  = 232;
  ram[69]  = 232;
  ram[70]  = 232;
  ram[71]  = 232;
  ram[72]  = 232;
  ram[73]  = 232;
  ram[74]  = 232;
  ram[75]  = 232;
  ram[76]  = 232;
  ram[77]  = 255;
  ram[78]  = 255;
  ram[79]  = 255;
  ram[80]  = 255;
  ram[81]  = 255;
  ram[82]  = 232;
  ram[83]  = 232;
  ram[84]  = 232;
  ram[85]  = 232;
  ram[86]  = 232;
  ram[87]  = 232;
  ram[88]  = 232;
  ram[89]  = 232;
  ram[90]  = 232;
  ram[91]  = 232;
  ram[92]  = 232;
  ram[93]  = 232;
  ram[94]  = 232;
  ram[95]  = 232;
  ram[96]  = 232;
  ram[97]  = 255;
  ram[98]  = 255;
  ram[99]  = 255;
  ram[100]  = 255;
  ram[101]  = 232;
  ram[102]  = 232;
  ram[103]  = 232;
  ram[104]  = 232;
  ram[105]  = 232;
  ram[106]  = 232;
  ram[107]  = 232;
  ram[108]  = 255;
  ram[109]  = 255;
  ram[110]  = 255;
  ram[111]  = 232;
  ram[112]  = 232;
  ram[113]  = 232;
  ram[114]  = 232;
  ram[115]  = 232;
  ram[116]  = 232;
  ram[117]  = 232;
  ram[118]  = 255;
  ram[119]  = 255;
  ram[120]  = 255;
  ram[121]  = 232;
  ram[122]  = 232;
  ram[123]  = 232;
  ram[124]  = 232;
  ram[125]  = 232;
  ram[126]  = 255;
  ram[127]  = 255;
  ram[128]  = 255;
  ram[129]  = 255;
  ram[130]  = 255;
  ram[131]  = 255;
  ram[132]  = 255;
  ram[133]  = 232;
  ram[134]  = 232;
  ram[135]  = 232;
  ram[136]  = 232;
  ram[137]  = 232;
  ram[138]  = 255;
  ram[139]  = 255;
  ram[140]  = 232;
  ram[141]  = 232;
  ram[142]  = 232;
  ram[143]  = 232;
  ram[144]  = 232;
  ram[145]  = 232;
  ram[146]  = 255;
  ram[147]  = 255;
  ram[148]  = 255;
  ram[149]  = 255;
  ram[150]  = 255;
  ram[151]  = 255;
  ram[152]  = 255;
  ram[153]  = 232;
  ram[154]  = 232;
  ram[155]  = 232;
  ram[156]  = 232;
  ram[157]  = 232;
  ram[158]  = 232;
  ram[159]  = 255;
  ram[160]  = 232;
  ram[161]  = 232;
  ram[162]  = 232;
  ram[163]  = 232;
  ram[164]  = 232;
  ram[165]  = 255;
  ram[166]  = 255;
  ram[167]  = 255;
  ram[168]  = 255;
  ram[169]  = 255;
  ram[170]  = 255;
  ram[171]  = 255;
  ram[172]  = 255;
  ram[173]  = 255;
  ram[174]  = 232;
  ram[175]  = 232;
  ram[176]  = 232;
  ram[177]  = 232;
  ram[178]  = 232;
  ram[179]  = 255;
  ram[180]  = 232;
  ram[181]  = 232;
  ram[182]  = 232;
  ram[183]  = 232;
  ram[184]  = 232;
  ram[185]  = 255;
  ram[186]  = 255;
  ram[187]  = 255;
  ram[188]  = 255;
  ram[189]  = 255;
  ram[190]  = 255;
  ram[191]  = 255;
  ram[192]  = 255;
  ram[193]  = 255;
  ram[194]  = 232;
  ram[195]  = 232;
  ram[196]  = 232;
  ram[197]  = 232;
  ram[198]  = 232;
  ram[199]  = 255;
  ram[200]  = 232;
  ram[201]  = 232;
  ram[202]  = 232;
  ram[203]  = 232;
  ram[204]  = 232;
  ram[205]  = 255;
  ram[206]  = 255;
  ram[207]  = 255;
  ram[208]  = 255;
  ram[209]  = 255;
  ram[210]  = 255;
  ram[211]  = 255;
  ram[212]  = 255;
  ram[213]  = 255;
  ram[214]  = 232;
  ram[215]  = 232;
  ram[216]  = 232;
  ram[217]  = 232;
  ram[218]  = 232;
  ram[219]  = 255;
  ram[220]  = 232;
  ram[221]  = 232;
  ram[222]  = 232;
  ram[223]  = 232;
  ram[224]  = 232;
  ram[225]  = 255;
  ram[226]  = 255;
  ram[227]  = 255;
  ram[228]  = 255;
  ram[229]  = 255;
  ram[230]  = 255;
  ram[231]  = 255;
  ram[232]  = 255;
  ram[233]  = 255;
  ram[234]  = 232;
  ram[235]  = 232;
  ram[236]  = 232;
  ram[237]  = 232;
  ram[238]  = 232;
  ram[239]  = 255;
  ram[240]  = 232;
  ram[241]  = 232;
  ram[242]  = 232;
  ram[243]  = 232;
  ram[244]  = 232;
  ram[245]  = 232;
  ram[246]  = 255;
  ram[247]  = 255;
  ram[248]  = 255;
  ram[249]  = 255;
  ram[250]  = 255;
  ram[251]  = 255;
  ram[252]  = 255;
  ram[253]  = 232;
  ram[254]  = 232;
  ram[255]  = 232;
  ram[256]  = 232;
  ram[257]  = 232;
  ram[258]  = 232;
  ram[259]  = 255;
  ram[260]  = 255;
  ram[261]  = 232;
  ram[262]  = 232;
  ram[263]  = 232;
  ram[264]  = 232;
  ram[265]  = 232;
  ram[266]  = 255;
  ram[267]  = 255;
  ram[268]  = 255;
  ram[269]  = 255;
  ram[270]  = 255;
  ram[271]  = 255;
  ram[272]  = 255;
  ram[273]  = 232;
  ram[274]  = 232;
  ram[275]  = 232;
  ram[276]  = 232;
  ram[277]  = 232;
  ram[278]  = 255;
  ram[279]  = 255;
  ram[280]  = 255;
  ram[281]  = 232;
  ram[282]  = 232;
  ram[283]  = 232;
  ram[284]  = 232;
  ram[285]  = 232;
  ram[286]  = 232;
  ram[287]  = 232;
  ram[288]  = 255;
  ram[289]  = 255;
  ram[290]  = 255;
  ram[291]  = 232;
  ram[292]  = 232;
  ram[293]  = 232;
  ram[294]  = 232;
  ram[295]  = 232;
  ram[296]  = 232;
  ram[297]  = 232;
  ram[298]  = 255;
  ram[299]  = 255;
  ram[300]  = 255;
  ram[301]  = 255;
  ram[302]  = 232;
  ram[303]  = 232;
  ram[304]  = 232;
  ram[305]  = 232;
  ram[306]  = 232;
  ram[307]  = 232;
  ram[308]  = 232;
  ram[309]  = 232;
  ram[310]  = 232;
  ram[311]  = 232;
  ram[312]  = 232;
  ram[313]  = 232;
  ram[314]  = 232;
  ram[315]  = 232;
  ram[316]  = 232;
  ram[317]  = 255;
  ram[318]  = 255;
  ram[319]  = 255;
  ram[320]  = 255;
  ram[321]  = 255;
  ram[322]  = 232;
  ram[323]  = 232;
  ram[324]  = 232;
  ram[325]  = 232;
  ram[326]  = 232;
  ram[327]  = 232;
  ram[328]  = 232;
  ram[329]  = 232;
  ram[330]  = 232;
  ram[331]  = 232;
  ram[332]  = 232;
  ram[333]  = 232;
  ram[334]  = 232;
  ram[335]  = 232;
  ram[336]  = 232;
  ram[337]  = 255;
  ram[338]  = 255;
  ram[339]  = 255;
  ram[340]  = 255;
  ram[341]  = 255;
  ram[342]  = 255;
  ram[343]  = 232;
  ram[344]  = 232;
  ram[345]  = 232;
  ram[346]  = 232;
  ram[347]  = 232;
  ram[348]  = 232;
  ram[349]  = 232;
  ram[350]  = 232;
  ram[351]  = 232;
  ram[352]  = 232;
  ram[353]  = 232;
  ram[354]  = 232;
  ram[355]  = 232;
  ram[356]  = 255;
  ram[357]  = 255;
  ram[358]  = 255;
  ram[359]  = 255;
  ram[360]  = 255;
  ram[361]  = 255;
  ram[362]  = 255;
  ram[363]  = 255;
  ram[364]  = 255;
  ram[365]  = 232;
  ram[366]  = 232;
  ram[367]  = 232;
  ram[368]  = 232;
  ram[369]  = 232;
  ram[370]  = 232;
  ram[371]  = 232;
  ram[372]  = 232;
  ram[373]  = 232;
  ram[374]  = 255;
  ram[375]  = 255;
  ram[376]  = 255;
  ram[377]  = 255;
  ram[378]  = 255;
  ram[379]  = 255;
  ram[380]  = 255;
  ram[381]  = 255;
  ram[382]  = 255;
  ram[383]  = 255;
  ram[384]  = 255;
  ram[385]  = 255;
  ram[386]  = 255;
  ram[387]  = 232;
  ram[388]  = 232;
  ram[389]  = 232;
  ram[390]  = 232;
  ram[391]  = 232;
  ram[392]  = 255;
  ram[393]  = 255;
  ram[394]  = 255;
  ram[395]  = 255;
  ram[396]  = 255;
  ram[397]  = 255;
  ram[398]  = 255;
  ram[399]  = 255;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
