module rom_man_g(clock, address, q);        // ROM-stored RGB bitmap for player(man)
input clock;
output [7:0] q;
input [8:0] address;
reg [7:0] dout;
reg [7:0] ram [511:0];
assign q = dout;

initial begin
  ram[0]  = 74;
  ram[1]  = 72;
  ram[2]  = 72;
  ram[3]  = 75;
  ram[4]  = 72;
  ram[5]  = 65;
  ram[6]  = 65;
  ram[7]  = 64;
  ram[8]  = 76;
  ram[9]  = 92;
  ram[10]  = 80;
  ram[11]  = 67;
  ram[12]  = 65;
  ram[13]  = 66;
  ram[14]  = 71;
  ram[15]  = 72;
  ram[16]  = 71;
  ram[17]  = 72;
  ram[18]  = 68;
  ram[19]  = 187;
  ram[20]  = 74;
  ram[21]  = 75;
  ram[22]  = 73;
  ram[23]  = 64;
  ram[24]  = 80;
  ram[25]  = 112;
  ram[26]  = 133;
  ram[27]  = 156;
  ram[28]  = 181;
  ram[29]  = 209;
  ram[30]  = 193;
  ram[31]  = 162;
  ram[32]  = 143;
  ram[33]  = 120;
  ram[34]  = 93;
  ram[35]  = 66;
  ram[36]  = 74;
  ram[37]  = 76;
  ram[38]  = 69;
  ram[39]  = 162;
  ram[40]  = 75;
  ram[41]  = 75;
  ram[42]  = 67;
  ram[43]  = 84;
  ram[44]  = 166;
  ram[45]  = 212;
  ram[46]  = 211;
  ram[47]  = 210;
  ram[48]  = 212;
  ram[49]  = 213;
  ram[50]  = 214;
  ram[51]  = 210;
  ram[52]  = 209;
  ram[53]  = 210;
  ram[54]  = 188;
  ram[55]  = 108;
  ram[56]  = 63;
  ram[57]  = 71;
  ram[58]  = 70;
  ram[59]  = 160;
  ram[60]  = 72;
  ram[61]  = 66;
  ram[62]  = 89;
  ram[63]  = 179;
  ram[64]  = 209;
  ram[65]  = 206;
  ram[66]  = 203;
  ram[67]  = 202;
  ram[68]  = 209;
  ram[69]  = 212;
  ram[70]  = 210;
  ram[71]  = 203;
  ram[72]  = 202;
  ram[73]  = 204;
  ram[74]  = 209;
  ram[75]  = 202;
  ram[76]  = 121;
  ram[77]  = 67;
  ram[78]  = 68;
  ram[79]  = 161;
  ram[80]  = 70;
  ram[81]  = 72;
  ram[82]  = 165;
  ram[83]  = 213;
  ram[84]  = 205;
  ram[85]  = 202;
  ram[86]  = 200;
  ram[87]  = 203;
  ram[88]  = 210;
  ram[89]  = 212;
  ram[90]  = 211;
  ram[91]  = 204;
  ram[92]  = 201;
  ram[93]  = 204;
  ram[94]  = 204;
  ram[95]  = 209;
  ram[96]  = 195;
  ram[97]  = 99;
  ram[98]  = 62;
  ram[99]  = 161;
  ram[100]  = 68;
  ram[101]  = 106;
  ram[102]  = 204;
  ram[103]  = 207;
  ram[104]  = 203;
  ram[105]  = 202;
  ram[106]  = 203;
  ram[107]  = 208;
  ram[108]  = 214;
  ram[109]  = 214;
  ram[110]  = 214;
  ram[111]  = 209;
  ram[112]  = 202;
  ram[113]  = 206;
  ram[114]  = 204;
  ram[115]  = 201;
  ram[116]  = 209;
  ram[117]  = 151;
  ram[118]  = 65;
  ram[119]  = 160;
  ram[120]  = 68;
  ram[121]  = 130;
  ram[122]  = 205;
  ram[123]  = 206;
  ram[124]  = 205;
  ram[125]  = 205;
  ram[126]  = 207;
  ram[127]  = 211;
  ram[128]  = 210;
  ram[129]  = 208;
  ram[130]  = 209;
  ram[131]  = 211;
  ram[132]  = 205;
  ram[133]  = 204;
  ram[134]  = 206;
  ram[135]  = 203;
  ram[136]  = 209;
  ram[137]  = 187;
  ram[138]  = 82;
  ram[139]  = 157;
  ram[140]  = 66;
  ram[141]  = 146;
  ram[142]  = 206;
  ram[143]  = 192;
  ram[144]  = 185;
  ram[145]  = 183;
  ram[146]  = 175;
  ram[147]  = 166;
  ram[148]  = 180;
  ram[149]  = 187;
  ram[150]  = 183;
  ram[151]  = 167;
  ram[152]  = 165;
  ram[153]  = 177;
  ram[154]  = 178;
  ram[155]  = 184;
  ram[156]  = 199;
  ram[157]  = 197;
  ram[158]  = 89;
  ram[159]  = 156;
  ram[160]  = 66;
  ram[161]  = 130;
  ram[162]  = 181;
  ram[163]  = 168;
  ram[164]  = 186;
  ram[165]  = 184;
  ram[166]  = 84;
  ram[167]  = 61;
  ram[168]  = 162;
  ram[169]  = 234;
  ram[170]  = 184;
  ram[171]  = 67;
  ram[172]  = 62;
  ram[173]  = 162;
  ram[174]  = 207;
  ram[175]  = 175;
  ram[176]  = 173;
  ram[177]  = 177;
  ram[178]  = 89;
  ram[179]  = 156;
  ram[180]  = 70;
  ram[181]  = 110;
  ram[182]  = 168;
  ram[183]  = 199;
  ram[184]  = 236;
  ram[185]  = 176;
  ram[186]  = 51;
  ram[187]  = 42;
  ram[188]  = 135;
  ram[189]  = 240;
  ram[190]  = 176;
  ram[191]  = 53;
  ram[192]  = 46;
  ram[193]  = 146;
  ram[194]  = 236;
  ram[195]  = 223;
  ram[196]  = 191;
  ram[197]  = 155;
  ram[198]  = 84;
  ram[199]  = 158;
  ram[200]  = 71;
  ram[201]  = 68;
  ram[202]  = 92;
  ram[203]  = 147;
  ram[204]  = 227;
  ram[205]  = 204;
  ram[206]  = 71;
  ram[207]  = 47;
  ram[208]  = 170;
  ram[209]  = 234;
  ram[210]  = 201;
  ram[211]  = 75;
  ram[212]  = 51;
  ram[213]  = 174;
  ram[214]  = 234;
  ram[215]  = 197;
  ram[216]  = 119;
  ram[217]  = 79;
  ram[218]  = 64;
  ram[219]  = 161;
  ram[220]  = 74;
  ram[221]  = 72;
  ram[222]  = 62;
  ram[223]  = 67;
  ram[224]  = 152;
  ram[225]  = 231;
  ram[226]  = 183;
  ram[227]  = 165;
  ram[228]  = 222;
  ram[229]  = 225;
  ram[230]  = 225;
  ram[231]  = 180;
  ram[232]  = 163;
  ram[233]  = 225;
  ram[234]  = 207;
  ram[235]  = 111;
  ram[236]  = 58;
  ram[237]  = 68;
  ram[238]  = 66;
  ram[239]  = 161;
  ram[240]  = 74;
  ram[241]  = 73;
  ram[242]  = 83;
  ram[243]  = 110;
  ram[244]  = 124;
  ram[245]  = 190;
  ram[246]  = 233;
  ram[247]  = 229;
  ram[248]  = 221;
  ram[249]  = 219;
  ram[250]  = 219;
  ram[251]  = 226;
  ram[252]  = 231;
  ram[253]  = 211;
  ram[254]  = 146;
  ram[255]  = 118;
  ram[256]  = 92;
  ram[257]  = 72;
  ram[258]  = 67;
  ram[259]  = 161;
  ram[260]  = 71;
  ram[261]  = 72;
  ram[262]  = 108;
  ram[263]  = 132;
  ram[264]  = 126;
  ram[265]  = 136;
  ram[266]  = 181;
  ram[267]  = 212;
  ram[268]  = 219;
  ram[269]  = 221;
  ram[270]  = 221;
  ram[271]  = 218;
  ram[272]  = 197;
  ram[273]  = 150;
  ram[274]  = 125;
  ram[275]  = 131;
  ram[276]  = 121;
  ram[277]  = 80;
  ram[278]  = 66;
  ram[279]  = 161;
  ram[280]  = 70;
  ram[281]  = 74;
  ram[282]  = 111;
  ram[283]  = 128;
  ram[284]  = 125;
  ram[285]  = 128;
  ram[286]  = 137;
  ram[287]  = 151;
  ram[288]  = 165;
  ram[289]  = 172;
  ram[290]  = 170;
  ram[291]  = 158;
  ram[292]  = 141;
  ram[293]  = 132;
  ram[294]  = 123;
  ram[295]  = 128;
  ram[296]  = 124;
  ram[297]  = 83;
  ram[298]  = 64;
  ram[299]  = 161;
  ram[300]  = 72;
  ram[301]  = 70;
  ram[302]  = 115;
  ram[303]  = 201;
  ram[304]  = 203;
  ram[305]  = 150;
  ram[306]  = 140;
  ram[307]  = 141;
  ram[308]  = 138;
  ram[309]  = 132;
  ram[310]  = 134;
  ram[311]  = 140;
  ram[312]  = 142;
  ram[313]  = 135;
  ram[314]  = 165;
  ram[315]  = 214;
  ram[316]  = 163;
  ram[317]  = 76;
  ram[318]  = 66;
  ram[319]  = 161;
  ram[320]  = 75;
  ram[321]  = 67;
  ram[322]  = 103;
  ram[323]  = 219;
  ram[324]  = 228;
  ram[325]  = 158;
  ram[326]  = 142;
  ram[327]  = 147;
  ram[328]  = 146;
  ram[329]  = 145;
  ram[330]  = 146;
  ram[331]  = 145;
  ram[332]  = 142;
  ram[333]  = 139;
  ram[334]  = 188;
  ram[335]  = 242;
  ram[336]  = 168;
  ram[337]  = 70;
  ram[338]  = 66;
  ram[339]  = 161;
  ram[340]  = 74;
  ram[341]  = 73;
  ram[342]  = 70;
  ram[343]  = 95;
  ram[344]  = 104;
  ram[345]  = 93;
  ram[346]  = 101;
  ram[347]  = 92;
  ram[348]  = 101;
  ram[349]  = 136;
  ram[350]  = 125;
  ram[351]  = 94;
  ram[352]  = 97;
  ram[353]  = 99;
  ram[354]  = 90;
  ram[355]  = 105;
  ram[356]  = 81;
  ram[357]  = 69;
  ram[358]  = 68;
  ram[359]  = 161;
  ram[360]  = 72;
  ram[361]  = 74;
  ram[362]  = 75;
  ram[363]  = 67;
  ram[364]  = 66;
  ram[365]  = 67;
  ram[366]  = 67;
  ram[367]  = 67;
  ram[368]  = 69;
  ram[369]  = 85;
  ram[370]  = 79;
  ram[371]  = 70;
  ram[372]  = 70;
  ram[373]  = 68;
  ram[374]  = 66;
  ram[375]  = 65;
  ram[376]  = 68;
  ram[377]  = 74;
  ram[378]  = 69;
  ram[379]  = 161;
  ram[380]  = 74;
  ram[381]  = 73;
  ram[382]  = 73;
  ram[383]  = 73;
  ram[384]  = 73;
  ram[385]  = 71;
  ram[386]  = 71;
  ram[387]  = 74;
  ram[388]  = 75;
  ram[389]  = 69;
  ram[390]  = 69;
  ram[391]  = 72;
  ram[392]  = 73;
  ram[393]  = 73;
  ram[394]  = 72;
  ram[395]  = 74;
  ram[396]  = 74;
  ram[397]  = 75;
  ram[398]  = 69;
  ram[399]  = 161;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
