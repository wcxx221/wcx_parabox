module rom_tui(clock, address, q);  // using rom to form display region 0
input clock;
output [7:0] q;
input [12:0] address;
reg [7:0] dout;
reg [7:0] ram [8191:0];
assign q = dout;

initial begin
  ram[0]  = 244;
  ram[1]  = 242;
  ram[2]  = 243;
  ram[3]  = 239;
  ram[4]  = 244;
  ram[5]  = 247;
  ram[6]  = 243;
  ram[7]  = 244;
  ram[8]  = 239;
  ram[9]  = 230;
  ram[10]  = 242;
  ram[11]  = 245;
  ram[12]  = 244;
  ram[13]  = 242;
  ram[14]  = 244;
  ram[15]  = 242;
  ram[16]  = 240;
  ram[17]  = 243;
  ram[18]  = 232;
  ram[19]  = 231;
  ram[20]  = 241;
  ram[21]  = 243;
  ram[22]  = 243;
  ram[23]  = 243;
  ram[24]  = 241;
  ram[25]  = 243;
  ram[26]  = 245;
  ram[27]  = 243;
  ram[28]  = 241;
  ram[29]  = 233;
  ram[30]  = 230;
  ram[31]  = 238;
  ram[32]  = 242;
  ram[33]  = 242;
  ram[34]  = 240;
  ram[35]  = 240;
  ram[36]  = 242;
  ram[37]  = 242;
  ram[38]  = 244;
  ram[39]  = 240;
  ram[40]  = 227;
  ram[41]  = 231;
  ram[42]  = 239;
  ram[43]  = 241;
  ram[44]  = 239;
  ram[45]  = 239;
  ram[46]  = 233;
  ram[47]  = 235;
  ram[48]  = 241;
  ram[49]  = 240;
  ram[50]  = 240;
  ram[51]  = 229;
  ram[52]  = 224;
  ram[53]  = 239;
  ram[54]  = 243;
  ram[55]  = 242;
  ram[56]  = 238;
  ram[57]  = 240;
  ram[58]  = 245;
  ram[59]  = 239;
  ram[60]  = 240;
  ram[61]  = 242;
  ram[62]  = 237;
  ram[63]  = 228;
  ram[64]  = 238;
  ram[65]  = 242;
  ram[66]  = 242;
  ram[67]  = 241;
  ram[68]  = 239;
  ram[69]  = 242;
  ram[70]  = 242;
  ram[71]  = 241;
  ram[72]  = 240;
  ram[73]  = 244;
  ram[74]  = 239;
  ram[75]  = 234;
  ram[76]  = 240;
  ram[77]  = 244;
  ram[78]  = 240;
  ram[79]  = 236;
  ram[80]  = 238;
  ram[81]  = 242;
  ram[82]  = 240;
  ram[83]  = 238;
  ram[84]  = 244;
  ram[85]  = 239;
  ram[86]  = 229;
  ram[87]  = 236;
  ram[88]  = 240;
  ram[89]  = 240;
  ram[90]  = 241;
  ram[91]  = 242;
  ram[92]  = 235;
  ram[93]  = 237;
  ram[94]  = 240;
  ram[95]  = 242;
  ram[96]  = 241;
  ram[97]  = 228;
  ram[98]  = 229;
  ram[99]  = 238;
  ram[100]  = 239;
  ram[101]  = 238;
  ram[102]  = 240;
  ram[103]  = 238;
  ram[104]  = 237;
  ram[105]  = 236;
  ram[106]  = 238;
  ram[107]  = 239;
  ram[108]  = 232;
  ram[109]  = 233;
  ram[110]  = 239;
  ram[111]  = 235;
  ram[112]  = 236;
  ram[113]  = 238;
  ram[114]  = 237;
  ram[115]  = 238;
  ram[116]  = 237;
  ram[117]  = 236;
  ram[118]  = 236;
  ram[119]  = 229;
  ram[120]  = 253;
  ram[121]  = 252;
  ram[122]  = 252;
  ram[123]  = 250;
  ram[124]  = 253;
  ram[125]  = 253;
  ram[126]  = 254;
  ram[127]  = 253;
  ram[128]  = 250;
  ram[129]  = 241;
  ram[130]  = 251;
  ram[131]  = 251;
  ram[132]  = 252;
  ram[133]  = 253;
  ram[134]  = 253;
  ram[135]  = 253;
  ram[136]  = 253;
  ram[137]  = 253;
  ram[138]  = 245;
  ram[139]  = 244;
  ram[140]  = 252;
  ram[141]  = 253;
  ram[142]  = 252;
  ram[143]  = 250;
  ram[144]  = 250;
  ram[145]  = 252;
  ram[146]  = 252;
  ram[147]  = 254;
  ram[148]  = 253;
  ram[149]  = 244;
  ram[150]  = 240;
  ram[151]  = 252;
  ram[152]  = 253;
  ram[153]  = 253;
  ram[154]  = 252;
  ram[155]  = 250;
  ram[156]  = 251;
  ram[157]  = 251;
  ram[158]  = 251;
  ram[159]  = 249;
  ram[160]  = 237;
  ram[161]  = 242;
  ram[162]  = 252;
  ram[163]  = 251;
  ram[164]  = 249;
  ram[165]  = 250;
  ram[166]  = 249;
  ram[167]  = 248;
  ram[168]  = 249;
  ram[169]  = 249;
  ram[170]  = 249;
  ram[171]  = 238;
  ram[172]  = 238;
  ram[173]  = 251;
  ram[174]  = 252;
  ram[175]  = 250;
  ram[176]  = 248;
  ram[177]  = 250;
  ram[178]  = 250;
  ram[179]  = 249;
  ram[180]  = 248;
  ram[181]  = 249;
  ram[182]  = 245;
  ram[183]  = 237;
  ram[184]  = 247;
  ram[185]  = 249;
  ram[186]  = 247;
  ram[187]  = 247;
  ram[188]  = 248;
  ram[189]  = 249;
  ram[190]  = 246;
  ram[191]  = 245;
  ram[192]  = 247;
  ram[193]  = 246;
  ram[194]  = 243;
  ram[195]  = 239;
  ram[196]  = 248;
  ram[197]  = 248;
  ram[198]  = 244;
  ram[199]  = 242;
  ram[200]  = 245;
  ram[201]  = 244;
  ram[202]  = 244;
  ram[203]  = 245;
  ram[204]  = 247;
  ram[205]  = 245;
  ram[206]  = 239;
  ram[207]  = 246;
  ram[208]  = 247;
  ram[209]  = 248;
  ram[210]  = 249;
  ram[211]  = 248;
  ram[212]  = 248;
  ram[213]  = 248;
  ram[214]  = 249;
  ram[215]  = 250;
  ram[216]  = 249;
  ram[217]  = 238;
  ram[218]  = 238;
  ram[219]  = 249;
  ram[220]  = 248;
  ram[221]  = 248;
  ram[222]  = 250;
  ram[223]  = 250;
  ram[224]  = 250;
  ram[225]  = 249;
  ram[226]  = 250;
  ram[227]  = 251;
  ram[228]  = 243;
  ram[229]  = 242;
  ram[230]  = 249;
  ram[231]  = 250;
  ram[232]  = 250;
  ram[233]  = 248;
  ram[234]  = 250;
  ram[235]  = 252;
  ram[236]  = 251;
  ram[237]  = 249;
  ram[238]  = 248;
  ram[239]  = 241;
  ram[240]  = 252;
  ram[241]  = 251;
  ram[242]  = 251;
  ram[243]  = 251;
  ram[244]  = 251;
  ram[245]  = 252;
  ram[246]  = 252;
  ram[247]  = 252;
  ram[248]  = 248;
  ram[249]  = 243;
  ram[250]  = 252;
  ram[251]  = 253;
  ram[252]  = 253;
  ram[253]  = 252;
  ram[254]  = 252;
  ram[255]  = 253;
  ram[256]  = 252;
  ram[257]  = 254;
  ram[258]  = 245;
  ram[259]  = 244;
  ram[260]  = 254;
  ram[261]  = 252;
  ram[262]  = 251;
  ram[263]  = 251;
  ram[264]  = 253;
  ram[265]  = 250;
  ram[266]  = 250;
  ram[267]  = 253;
  ram[268]  = 251;
  ram[269]  = 243;
  ram[270]  = 241;
  ram[271]  = 251;
  ram[272]  = 252;
  ram[273]  = 253;
  ram[274]  = 253;
  ram[275]  = 252;
  ram[276]  = 253;
  ram[277]  = 252;
  ram[278]  = 252;
  ram[279]  = 251;
  ram[280]  = 239;
  ram[281]  = 247;
  ram[282]  = 255;
  ram[283]  = 253;
  ram[284]  = 250;
  ram[285]  = 250;
  ram[286]  = 252;
  ram[287]  = 253;
  ram[288]  = 252;
  ram[289]  = 252;
  ram[290]  = 252;
  ram[291]  = 241;
  ram[292]  = 244;
  ram[293]  = 255;
  ram[294]  = 253;
  ram[295]  = 251;
  ram[296]  = 251;
  ram[297]  = 254;
  ram[298]  = 252;
  ram[299]  = 251;
  ram[300]  = 250;
  ram[301]  = 252;
  ram[302]  = 249;
  ram[303]  = 242;
  ram[304]  = 250;
  ram[305]  = 253;
  ram[306]  = 252;
  ram[307]  = 253;
  ram[308]  = 254;
  ram[309]  = 251;
  ram[310]  = 249;
  ram[311]  = 253;
  ram[312]  = 253;
  ram[313]  = 253;
  ram[314]  = 250;
  ram[315]  = 244;
  ram[316]  = 252;
  ram[317]  = 252;
  ram[318]  = 251;
  ram[319]  = 253;
  ram[320]  = 253;
  ram[321]  = 251;
  ram[322]  = 251;
  ram[323]  = 253;
  ram[324]  = 254;
  ram[325]  = 249;
  ram[326]  = 243;
  ram[327]  = 252;
  ram[328]  = 252;
  ram[329]  = 253;
  ram[330]  = 252;
  ram[331]  = 253;
  ram[332]  = 252;
  ram[333]  = 252;
  ram[334]  = 253;
  ram[335]  = 253;
  ram[336]  = 252;
  ram[337]  = 242;
  ram[338]  = 240;
  ram[339]  = 252;
  ram[340]  = 251;
  ram[341]  = 251;
  ram[342]  = 252;
  ram[343]  = 253;
  ram[344]  = 253;
  ram[345]  = 252;
  ram[346]  = 251;
  ram[347]  = 253;
  ram[348]  = 247;
  ram[349]  = 245;
  ram[350]  = 252;
  ram[351]  = 252;
  ram[352]  = 252;
  ram[353]  = 251;
  ram[354]  = 253;
  ram[355]  = 252;
  ram[356]  = 253;
  ram[357]  = 252;
  ram[358]  = 251;
  ram[359]  = 246;
  ram[360]  = 252;
  ram[361]  = 250;
  ram[362]  = 251;
  ram[363]  = 250;
  ram[364]  = 251;
  ram[365]  = 251;
  ram[366]  = 251;
  ram[367]  = 251;
  ram[368]  = 249;
  ram[369]  = 243;
  ram[370]  = 251;
  ram[371]  = 253;
  ram[372]  = 253;
  ram[373]  = 252;
  ram[374]  = 252;
  ram[375]  = 253;
  ram[376]  = 253;
  ram[377]  = 253;
  ram[378]  = 246;
  ram[379]  = 245;
  ram[380]  = 253;
  ram[381]  = 252;
  ram[382]  = 251;
  ram[383]  = 252;
  ram[384]  = 252;
  ram[385]  = 252;
  ram[386]  = 252;
  ram[387]  = 252;
  ram[388]  = 251;
  ram[389]  = 243;
  ram[390]  = 241;
  ram[391]  = 251;
  ram[392]  = 252;
  ram[393]  = 252;
  ram[394]  = 252;
  ram[395]  = 253;
  ram[396]  = 253;
  ram[397]  = 252;
  ram[398]  = 251;
  ram[399]  = 252;
  ram[400]  = 239;
  ram[401]  = 247;
  ram[402]  = 252;
  ram[403]  = 251;
  ram[404]  = 250;
  ram[405]  = 250;
  ram[406]  = 252;
  ram[407]  = 252;
  ram[408]  = 250;
  ram[409]  = 252;
  ram[410]  = 253;
  ram[411]  = 244;
  ram[412]  = 242;
  ram[413]  = 253;
  ram[414]  = 252;
  ram[415]  = 250;
  ram[416]  = 250;
  ram[417]  = 252;
  ram[418]  = 251;
  ram[419]  = 249;
  ram[420]  = 250;
  ram[421]  = 251;
  ram[422]  = 249;
  ram[423]  = 241;
  ram[424]  = 255;
  ram[425]  = 255;
  ram[426]  = 255;
  ram[427]  = 252;
  ram[428]  = 251;
  ram[429]  = 250;
  ram[430]  = 249;
  ram[431]  = 251;
  ram[432]  = 252;
  ram[433]  = 253;
  ram[434]  = 249;
  ram[435]  = 243;
  ram[436]  = 251;
  ram[437]  = 250;
  ram[438]  = 250;
  ram[439]  = 251;
  ram[440]  = 251;
  ram[441]  = 249;
  ram[442]  = 248;
  ram[443]  = 253;
  ram[444]  = 253;
  ram[445]  = 248;
  ram[446]  = 240;
  ram[447]  = 251;
  ram[448]  = 252;
  ram[449]  = 252;
  ram[450]  = 252;
  ram[451]  = 253;
  ram[452]  = 251;
  ram[453]  = 251;
  ram[454]  = 252;
  ram[455]  = 252;
  ram[456]  = 252;
  ram[457]  = 243;
  ram[458]  = 243;
  ram[459]  = 252;
  ram[460]  = 253;
  ram[461]  = 251;
  ram[462]  = 251;
  ram[463]  = 252;
  ram[464]  = 252;
  ram[465]  = 252;
  ram[466]  = 251;
  ram[467]  = 253;
  ram[468]  = 245;
  ram[469]  = 244;
  ram[470]  = 251;
  ram[471]  = 250;
  ram[472]  = 250;
  ram[473]  = 250;
  ram[474]  = 252;
  ram[475]  = 252;
  ram[476]  = 252;
  ram[477]  = 249;
  ram[478]  = 250;
  ram[479]  = 246;
  ram[480]  = 251;
  ram[481]  = 251;
  ram[482]  = 251;
  ram[483]  = 250;
  ram[484]  = 250;
  ram[485]  = 250;
  ram[486]  = 250;
  ram[487]  = 251;
  ram[488]  = 248;
  ram[489]  = 239;
  ram[490]  = 251;
  ram[491]  = 252;
  ram[492]  = 253;
  ram[493]  = 253;
  ram[494]  = 252;
  ram[495]  = 252;
  ram[496]  = 253;
  ram[497]  = 253;
  ram[498]  = 245;
  ram[499]  = 245;
  ram[500]  = 253;
  ram[501]  = 253;
  ram[502]  = 252;
  ram[503]  = 252;
  ram[504]  = 255;
  ram[505]  = 255;
  ram[506]  = 255;
  ram[507]  = 252;
  ram[508]  = 252;
  ram[509]  = 246;
  ram[510]  = 241;
  ram[511]  = 251;
  ram[512]  = 253;
  ram[513]  = 252;
  ram[514]  = 251;
  ram[515]  = 252;
  ram[516]  = 253;
  ram[517]  = 252;
  ram[518]  = 252;
  ram[519]  = 252;
  ram[520]  = 238;
  ram[521]  = 246;
  ram[522]  = 251;
  ram[523]  = 250;
  ram[524]  = 251;
  ram[525]  = 251;
  ram[526]  = 252;
  ram[527]  = 251;
  ram[528]  = 253;
  ram[529]  = 253;
  ram[530]  = 253;
  ram[531]  = 255;
  ram[532]  = 255;
  ram[533]  = 255;
  ram[534]  = 252;
  ram[535]  = 251;
  ram[536]  = 251;
  ram[537]  = 251;
  ram[538]  = 251;
  ram[539]  = 252;
  ram[540]  = 251;
  ram[541]  = 250;
  ram[542]  = 248;
  ram[543]  = 250;
  ram[544]  = 174;
  ram[545]  = 114;
  ram[546]  = 191;
  ram[547]  = 252;
  ram[548]  = 253;
  ram[549]  = 250;
  ram[550]  = 251;
  ram[551]  = 252;
  ram[552]  = 252;
  ram[553]  = 253;
  ram[554]  = 248;
  ram[555]  = 242;
  ram[556]  = 249;
  ram[557]  = 250;
  ram[558]  = 249;
  ram[559]  = 250;
  ram[560]  = 250;
  ram[561]  = 249;
  ram[562]  = 249;
  ram[563]  = 252;
  ram[564]  = 251;
  ram[565]  = 249;
  ram[566]  = 241;
  ram[567]  = 251;
  ram[568]  = 252;
  ram[569]  = 252;
  ram[570]  = 252;
  ram[571]  = 253;
  ram[572]  = 252;
  ram[573]  = 252;
  ram[574]  = 253;
  ram[575]  = 253;
  ram[576]  = 253;
  ram[577]  = 244;
  ram[578]  = 243;
  ram[579]  = 253;
  ram[580]  = 253;
  ram[581]  = 252;
  ram[582]  = 252;
  ram[583]  = 252;
  ram[584]  = 252;
  ram[585]  = 253;
  ram[586]  = 253;
  ram[587]  = 254;
  ram[588]  = 245;
  ram[589]  = 243;
  ram[590]  = 251;
  ram[591]  = 249;
  ram[592]  = 251;
  ram[593]  = 250;
  ram[594]  = 251;
  ram[595]  = 252;
  ram[596]  = 252;
  ram[597]  = 251;
  ram[598]  = 251;
  ram[599]  = 248;
  ram[600]  = 250;
  ram[601]  = 251;
  ram[602]  = 251;
  ram[603]  = 251;
  ram[604]  = 249;
  ram[605]  = 251;
  ram[606]  = 251;
  ram[607]  = 254;
  ram[608]  = 249;
  ram[609]  = 239;
  ram[610]  = 251;
  ram[611]  = 253;
  ram[612]  = 253;
  ram[613]  = 255;
  ram[614]  = 253;
  ram[615]  = 252;
  ram[616]  = 253;
  ram[617]  = 253;
  ram[618]  = 245;
  ram[619]  = 246;
  ram[620]  = 252;
  ram[621]  = 253;
  ram[622]  = 253;
  ram[623]  = 255;
  ram[624]  = 212;
  ram[625]  = 181;
  ram[626]  = 255;
  ram[627]  = 254;
  ram[628]  = 253;
  ram[629]  = 245;
  ram[630]  = 242;
  ram[631]  = 252;
  ram[632]  = 252;
  ram[633]  = 253;
  ram[634]  = 252;
  ram[635]  = 252;
  ram[636]  = 252;
  ram[637]  = 252;
  ram[638]  = 253;
  ram[639]  = 252;
  ram[640]  = 239;
  ram[641]  = 246;
  ram[642]  = 251;
  ram[643]  = 250;
  ram[644]  = 252;
  ram[645]  = 252;
  ram[646]  = 250;
  ram[647]  = 251;
  ram[648]  = 252;
  ram[649]  = 253;
  ram[650]  = 255;
  ram[651]  = 180;
  ram[652]  = 164;
  ram[653]  = 244;
  ram[654]  = 255;
  ram[655]  = 252;
  ram[656]  = 252;
  ram[657]  = 252;
  ram[658]  = 251;
  ram[659]  = 253;
  ram[660]  = 251;
  ram[661]  = 251;
  ram[662]  = 254;
  ram[663]  = 243;
  ram[664]  = 30;
  ram[665]  = 0;
  ram[666]  = 0;
  ram[667]  = 171;
  ram[668]  = 255;
  ram[669]  = 253;
  ram[670]  = 252;
  ram[671]  = 253;
  ram[672]  = 253;
  ram[673]  = 254;
  ram[674]  = 249;
  ram[675]  = 242;
  ram[676]  = 250;
  ram[677]  = 250;
  ram[678]  = 249;
  ram[679]  = 251;
  ram[680]  = 251;
  ram[681]  = 249;
  ram[682]  = 251;
  ram[683]  = 252;
  ram[684]  = 252;
  ram[685]  = 248;
  ram[686]  = 242;
  ram[687]  = 251;
  ram[688]  = 252;
  ram[689]  = 251;
  ram[690]  = 252;
  ram[691]  = 252;
  ram[692]  = 253;
  ram[693]  = 252;
  ram[694]  = 252;
  ram[695]  = 253;
  ram[696]  = 254;
  ram[697]  = 246;
  ram[698]  = 248;
  ram[699]  = 255;
  ram[700]  = 255;
  ram[701]  = 255;
  ram[702]  = 255;
  ram[703]  = 255;
  ram[704]  = 254;
  ram[705]  = 252;
  ram[706]  = 253;
  ram[707]  = 254;
  ram[708]  = 245;
  ram[709]  = 244;
  ram[710]  = 249;
  ram[711]  = 248;
  ram[712]  = 252;
  ram[713]  = 251;
  ram[714]  = 250;
  ram[715]  = 252;
  ram[716]  = 252;
  ram[717]  = 252;
  ram[718]  = 252;
  ram[719]  = 248;
  ram[720]  = 251;
  ram[721]  = 252;
  ram[722]  = 252;
  ram[723]  = 250;
  ram[724]  = 250;
  ram[725]  = 251;
  ram[726]  = 252;
  ram[727]  = 253;
  ram[728]  = 251;
  ram[729]  = 240;
  ram[730]  = 251;
  ram[731]  = 253;
  ram[732]  = 255;
  ram[733]  = 244;
  ram[734]  = 255;
  ram[735]  = 255;
  ram[736]  = 253;
  ram[737]  = 253;
  ram[738]  = 246;
  ram[739]  = 246;
  ram[740]  = 252;
  ram[741]  = 252;
  ram[742]  = 255;
  ram[743]  = 227;
  ram[744]  = 26;
  ram[745]  = 0;
  ram[746]  = 92;
  ram[747]  = 250;
  ram[748]  = 254;
  ram[749]  = 255;
  ram[750]  = 255;
  ram[751]  = 255;
  ram[752]  = 253;
  ram[753]  = 252;
  ram[754]  = 253;
  ram[755]  = 252;
  ram[756]  = 251;
  ram[757]  = 252;
  ram[758]  = 253;
  ram[759]  = 252;
  ram[760]  = 240;
  ram[761]  = 246;
  ram[762]  = 252;
  ram[763]  = 250;
  ram[764]  = 253;
  ram[765]  = 252;
  ram[766]  = 250;
  ram[767]  = 251;
  ram[768]  = 251;
  ram[769]  = 255;
  ram[770]  = 228;
  ram[771]  = 9;
  ram[772]  = 0;
  ram[773]  = 51;
  ram[774]  = 232;
  ram[775]  = 255;
  ram[776]  = 253;
  ram[777]  = 251;
  ram[778]  = 253;
  ram[779]  = 254;
  ram[780]  = 253;
  ram[781]  = 251;
  ram[782]  = 255;
  ram[783]  = 165;
  ram[784]  = 1;
  ram[785]  = 0;
  ram[786]  = 0;
  ram[787]  = 129;
  ram[788]  = 255;
  ram[789]  = 255;
  ram[790]  = 255;
  ram[791]  = 255;
  ram[792]  = 255;
  ram[793]  = 255;
  ram[794]  = 255;
  ram[795]  = 243;
  ram[796]  = 249;
  ram[797]  = 251;
  ram[798]  = 250;
  ram[799]  = 250;
  ram[800]  = 251;
  ram[801]  = 250;
  ram[802]  = 251;
  ram[803]  = 252;
  ram[804]  = 253;
  ram[805]  = 249;
  ram[806]  = 243;
  ram[807]  = 251;
  ram[808]  = 251;
  ram[809]  = 251;
  ram[810]  = 253;
  ram[811]  = 255;
  ram[812]  = 255;
  ram[813]  = 255;
  ram[814]  = 255;
  ram[815]  = 255;
  ram[816]  = 255;
  ram[817]  = 255;
  ram[818]  = 249;
  ram[819]  = 226;
  ram[820]  = 230;
  ram[821]  = 219;
  ram[822]  = 219;
  ram[823]  = 204;
  ram[824]  = 255;
  ram[825]  = 255;
  ram[826]  = 253;
  ram[827]  = 253;
  ram[828]  = 248;
  ram[829]  = 247;
  ram[830]  = 250;
  ram[831]  = 249;
  ram[832]  = 249;
  ram[833]  = 250;
  ram[834]  = 249;
  ram[835]  = 252;
  ram[836]  = 251;
  ram[837]  = 253;
  ram[838]  = 252;
  ram[839]  = 245;
  ram[840]  = 251;
  ram[841]  = 252;
  ram[842]  = 251;
  ram[843]  = 250;
  ram[844]  = 250;
  ram[845]  = 251;
  ram[846]  = 252;
  ram[847]  = 252;
  ram[848]  = 249;
  ram[849]  = 240;
  ram[850]  = 250;
  ram[851]  = 255;
  ram[852]  = 190;
  ram[853]  = 59;
  ram[854]  = 71;
  ram[855]  = 212;
  ram[856]  = 255;
  ram[857]  = 253;
  ram[858]  = 246;
  ram[859]  = 247;
  ram[860]  = 254;
  ram[861]  = 252;
  ram[862]  = 255;
  ram[863]  = 128;
  ram[864]  = 0;
  ram[865]  = 0;
  ram[866]  = 34;
  ram[867]  = 249;
  ram[868]  = 255;
  ram[869]  = 218;
  ram[870]  = 134;
  ram[871]  = 221;
  ram[872]  = 255;
  ram[873]  = 253;
  ram[874]  = 252;
  ram[875]  = 252;
  ram[876]  = 252;
  ram[877]  = 253;
  ram[878]  = 253;
  ram[879]  = 252;
  ram[880]  = 240;
  ram[881]  = 246;
  ram[882]  = 253;
  ram[883]  = 252;
  ram[884]  = 251;
  ram[885]  = 251;
  ram[886]  = 251;
  ram[887]  = 251;
  ram[888]  = 251;
  ram[889]  = 255;
  ram[890]  = 137;
  ram[891]  = 0;
  ram[892]  = 0;
  ram[893]  = 0;
  ram[894]  = 182;
  ram[895]  = 255;
  ram[896]  = 255;
  ram[897]  = 255;
  ram[898]  = 255;
  ram[899]  = 255;
  ram[900]  = 255;
  ram[901]  = 254;
  ram[902]  = 255;
  ram[903]  = 76;
  ram[904]  = 0;
  ram[905]  = 0;
  ram[906]  = 0;
  ram[907]  = 141;
  ram[908]  = 210;
  ram[909]  = 167;
  ram[910]  = 139;
  ram[911]  = 115;
  ram[912]  = 94;
  ram[913]  = 94;
  ram[914]  = 210;
  ram[915]  = 253;
  ram[916]  = 250;
  ram[917]  = 252;
  ram[918]  = 251;
  ram[919]  = 250;
  ram[920]  = 250;
  ram[921]  = 251;
  ram[922]  = 252;
  ram[923]  = 252;
  ram[924]  = 253;
  ram[925]  = 248;
  ram[926]  = 242;
  ram[927]  = 252;
  ram[928]  = 255;
  ram[929]  = 255;
  ram[930]  = 255;
  ram[931]  = 245;
  ram[932]  = 222;
  ram[933]  = 201;
  ram[934]  = 151;
  ram[935]  = 126;
  ram[936]  = 83;
  ram[937]  = 74;
  ram[938]  = 50;
  ram[939]  = 15;
  ram[940]  = 19;
  ram[941]  = 11;
  ram[942]  = 15;
  ram[943]  = 4;
  ram[944]  = 90;
  ram[945]  = 224;
  ram[946]  = 255;
  ram[947]  = 254;
  ram[948]  = 246;
  ram[949]  = 242;
  ram[950]  = 251;
  ram[951]  = 250;
  ram[952]  = 249;
  ram[953]  = 250;
  ram[954]  = 249;
  ram[955]  = 250;
  ram[956]  = 251;
  ram[957]  = 252;
  ram[958]  = 250;
  ram[959]  = 246;
  ram[960]  = 252;
  ram[961]  = 252;
  ram[962]  = 252;
  ram[963]  = 250;
  ram[964]  = 250;
  ram[965]  = 252;
  ram[966]  = 253;
  ram[967]  = 252;
  ram[968]  = 249;
  ram[969]  = 241;
  ram[970]  = 253;
  ram[971]  = 255;
  ram[972]  = 70;
  ram[973]  = 0;
  ram[974]  = 0;
  ram[975]  = 119;
  ram[976]  = 255;
  ram[977]  = 254;
  ram[978]  = 245;
  ram[979]  = 247;
  ram[980]  = 254;
  ram[981]  = 255;
  ram[982]  = 245;
  ram[983]  = 35;
  ram[984]  = 0;
  ram[985]  = 0;
  ram[986]  = 92;
  ram[987]  = 255;
  ram[988]  = 252;
  ram[989]  = 51;
  ram[990]  = 0;
  ram[991]  = 19;
  ram[992]  = 166;
  ram[993]  = 255;
  ram[994]  = 253;
  ram[995]  = 251;
  ram[996]  = 252;
  ram[997]  = 253;
  ram[998]  = 253;
  ram[999]  = 253;
  ram[1000]  = 240;
  ram[1001]  = 247;
  ram[1002]  = 253;
  ram[1003]  = 252;
  ram[1004]  = 251;
  ram[1005]  = 251;
  ram[1006]  = 252;
  ram[1007]  = 251;
  ram[1008]  = 254;
  ram[1009]  = 248;
  ram[1010]  = 37;
  ram[1011]  = 0;
  ram[1012]  = 0;
  ram[1013]  = 12;
  ram[1014]  = 193;
  ram[1015]  = 205;
  ram[1016]  = 161;
  ram[1017]  = 139;
  ram[1018]  = 100;
  ram[1019]  = 86;
  ram[1020]  = 181;
  ram[1021]  = 255;
  ram[1022]  = 217;
  ram[1023]  = 9;
  ram[1024]  = 0;
  ram[1025]  = 0;
  ram[1026]  = 0;
  ram[1027]  = 12;
  ram[1028]  = 2;
  ram[1029]  = 0;
  ram[1030]  = 0;
  ram[1031]  = 0;
  ram[1032]  = 0;
  ram[1033]  = 0;
  ram[1034]  = 36;
  ram[1035]  = 239;
  ram[1036]  = 254;
  ram[1037]  = 253;
  ram[1038]  = 251;
  ram[1039]  = 251;
  ram[1040]  = 251;
  ram[1041]  = 253;
  ram[1042]  = 252;
  ram[1043]  = 252;
  ram[1044]  = 253;
  ram[1045]  = 248;
  ram[1046]  = 243;
  ram[1047]  = 253;
  ram[1048]  = 241;
  ram[1049]  = 154;
  ram[1050]  = 90;
  ram[1051]  = 37;
  ram[1052]  = 12;
  ram[1053]  = 1;
  ram[1054]  = 0;
  ram[1055]  = 0;
  ram[1056]  = 0;
  ram[1057]  = 0;
  ram[1058]  = 0;
  ram[1059]  = 0;
  ram[1060]  = 0;
  ram[1061]  = 0;
  ram[1062]  = 0;
  ram[1063]  = 0;
  ram[1064]  = 0;
  ram[1065]  = 36;
  ram[1066]  = 200;
  ram[1067]  = 255;
  ram[1068]  = 247;
  ram[1069]  = 243;
  ram[1070]  = 253;
  ram[1071]  = 252;
  ram[1072]  = 251;
  ram[1073]  = 250;
  ram[1074]  = 250;
  ram[1075]  = 249;
  ram[1076]  = 250;
  ram[1077]  = 250;
  ram[1078]  = 251;
  ram[1079]  = 246;
  ram[1080]  = 253;
  ram[1081]  = 251;
  ram[1082]  = 251;
  ram[1083]  = 251;
  ram[1084]  = 251;
  ram[1085]  = 252;
  ram[1086]  = 253;
  ram[1087]  = 253;
  ram[1088]  = 250;
  ram[1089]  = 242;
  ram[1090]  = 254;
  ram[1091]  = 254;
  ram[1092]  = 60;
  ram[1093]  = 0;
  ram[1094]  = 0;
  ram[1095]  = 72;
  ram[1096]  = 255;
  ram[1097]  = 255;
  ram[1098]  = 244;
  ram[1099]  = 247;
  ram[1100]  = 253;
  ram[1101]  = 255;
  ram[1102]  = 162;
  ram[1103]  = 0;
  ram[1104]  = 0;
  ram[1105]  = 0;
  ram[1106]  = 142;
  ram[1107]  = 255;
  ram[1108]  = 251;
  ram[1109]  = 61;
  ram[1110]  = 0;
  ram[1111]  = 0;
  ram[1112]  = 3;
  ram[1113]  = 177;
  ram[1114]  = 255;
  ram[1115]  = 252;
  ram[1116]  = 252;
  ram[1117]  = 253;
  ram[1118]  = 253;
  ram[1119]  = 253;
  ram[1120]  = 238;
  ram[1121]  = 246;
  ram[1122]  = 253;
  ram[1123]  = 252;
  ram[1124]  = 252;
  ram[1125]  = 252;
  ram[1126]  = 253;
  ram[1127]  = 252;
  ram[1128]  = 255;
  ram[1129]  = 170;
  ram[1130]  = 0;
  ram[1131]  = 0;
  ram[1132]  = 0;
  ram[1133]  = 6;
  ram[1134]  = 18;
  ram[1135]  = 0;
  ram[1136]  = 0;
  ram[1137]  = 0;
  ram[1138]  = 0;
  ram[1139]  = 0;
  ram[1140]  = 0;
  ram[1141]  = 214;
  ram[1142]  = 141;
  ram[1143]  = 0;
  ram[1144]  = 0;
  ram[1145]  = 0;
  ram[1146]  = 0;
  ram[1147]  = 0;
  ram[1148]  = 0;
  ram[1149]  = 0;
  ram[1150]  = 0;
  ram[1151]  = 0;
  ram[1152]  = 0;
  ram[1153]  = 0;
  ram[1154]  = 75;
  ram[1155]  = 236;
  ram[1156]  = 254;
  ram[1157]  = 253;
  ram[1158]  = 252;
  ram[1159]  = 251;
  ram[1160]  = 252;
  ram[1161]  = 252;
  ram[1162]  = 252;
  ram[1163]  = 252;
  ram[1164]  = 253;
  ram[1165]  = 249;
  ram[1166]  = 244;
  ram[1167]  = 255;
  ram[1168]  = 176;
  ram[1169]  = 0;
  ram[1170]  = 0;
  ram[1171]  = 0;
  ram[1172]  = 0;
  ram[1173]  = 0;
  ram[1174]  = 0;
  ram[1175]  = 0;
  ram[1176]  = 0;
  ram[1177]  = 0;
  ram[1178]  = 0;
  ram[1179]  = 0;
  ram[1180]  = 0;
  ram[1181]  = 0;
  ram[1182]  = 0;
  ram[1183]  = 0;
  ram[1184]  = 0;
  ram[1185]  = 0;
  ram[1186]  = 116;
  ram[1187]  = 255;
  ram[1188]  = 246;
  ram[1189]  = 246;
  ram[1190]  = 255;
  ram[1191]  = 252;
  ram[1192]  = 251;
  ram[1193]  = 250;
  ram[1194]  = 248;
  ram[1195]  = 249;
  ram[1196]  = 249;
  ram[1197]  = 249;
  ram[1198]  = 252;
  ram[1199]  = 247;
  ram[1200]  = 253;
  ram[1201]  = 252;
  ram[1202]  = 252;
  ram[1203]  = 251;
  ram[1204]  = 252;
  ram[1205]  = 253;
  ram[1206]  = 252;
  ram[1207]  = 253;
  ram[1208]  = 251;
  ram[1209]  = 244;
  ram[1210]  = 254;
  ram[1211]  = 255;
  ram[1212]  = 65;
  ram[1213]  = 0;
  ram[1214]  = 0;
  ram[1215]  = 47;
  ram[1216]  = 252;
  ram[1217]  = 255;
  ram[1218]  = 244;
  ram[1219]  = 247;
  ram[1220]  = 255;
  ram[1221]  = 244;
  ram[1222]  = 45;
  ram[1223]  = 0;
  ram[1224]  = 0;
  ram[1225]  = 24;
  ram[1226]  = 236;
  ram[1227]  = 255;
  ram[1228]  = 255;
  ram[1229]  = 175;
  ram[1230]  = 0;
  ram[1231]  = 0;
  ram[1232]  = 0;
  ram[1233]  = 11;
  ram[1234]  = 223;
  ram[1235]  = 255;
  ram[1236]  = 252;
  ram[1237]  = 252;
  ram[1238]  = 253;
  ram[1239]  = 253;
  ram[1240]  = 242;
  ram[1241]  = 247;
  ram[1242]  = 253;
  ram[1243]  = 251;
  ram[1244]  = 252;
  ram[1245]  = 253;
  ram[1246]  = 252;
  ram[1247]  = 255;
  ram[1248]  = 248;
  ram[1249]  = 37;
  ram[1250]  = 0;
  ram[1251]  = 0;
  ram[1252]  = 0;
  ram[1253]  = 0;
  ram[1254]  = 0;
  ram[1255]  = 0;
  ram[1256]  = 0;
  ram[1257]  = 0;
  ram[1258]  = 0;
  ram[1259]  = 0;
  ram[1260]  = 64;
  ram[1261]  = 232;
  ram[1262]  = 47;
  ram[1263]  = 0;
  ram[1264]  = 0;
  ram[1265]  = 5;
  ram[1266]  = 19;
  ram[1267]  = 0;
  ram[1268]  = 0;
  ram[1269]  = 49;
  ram[1270]  = 81;
  ram[1271]  = 107;
  ram[1272]  = 127;
  ram[1273]  = 168;
  ram[1274]  = 247;
  ram[1275]  = 248;
  ram[1276]  = 250;
  ram[1277]  = 253;
  ram[1278]  = 252;
  ram[1279]  = 251;
  ram[1280]  = 252;
  ram[1281]  = 252;
  ram[1282]  = 252;
  ram[1283]  = 252;
  ram[1284]  = 253;
  ram[1285]  = 249;
  ram[1286]  = 240;
  ram[1287]  = 255;
  ram[1288]  = 206;
  ram[1289]  = 14;
  ram[1290]  = 0;
  ram[1291]  = 0;
  ram[1292]  = 0;
  ram[1293]  = 0;
  ram[1294]  = 0;
  ram[1295]  = 0;
  ram[1296]  = 0;
  ram[1297]  = 11;
  ram[1298]  = 25;
  ram[1299]  = 65;
  ram[1300]  = 79;
  ram[1301]  = 0;
  ram[1302]  = 0;
  ram[1303]  = 0;
  ram[1304]  = 0;
  ram[1305]  = 0;
  ram[1306]  = 163;
  ram[1307]  = 255;
  ram[1308]  = 245;
  ram[1309]  = 246;
  ram[1310]  = 253;
  ram[1311]  = 250;
  ram[1312]  = 250;
  ram[1313]  = 251;
  ram[1314]  = 250;
  ram[1315]  = 250;
  ram[1316]  = 250;
  ram[1317]  = 250;
  ram[1318]  = 253;
  ram[1319]  = 244;
  ram[1320]  = 253;
  ram[1321]  = 252;
  ram[1322]  = 253;
  ram[1323]  = 253;
  ram[1324]  = 253;
  ram[1325]  = 253;
  ram[1326]  = 253;
  ram[1327]  = 254;
  ram[1328]  = 252;
  ram[1329]  = 246;
  ram[1330]  = 254;
  ram[1331]  = 255;
  ram[1332]  = 93;
  ram[1333]  = 0;
  ram[1334]  = 0;
  ram[1335]  = 26;
  ram[1336]  = 246;
  ram[1337]  = 255;
  ram[1338]  = 250;
  ram[1339]  = 249;
  ram[1340]  = 255;
  ram[1341]  = 176;
  ram[1342]  = 0;
  ram[1343]  = 0;
  ram[1344]  = 0;
  ram[1345]  = 125;
  ram[1346]  = 255;
  ram[1347]  = 255;
  ram[1348]  = 255;
  ram[1349]  = 251;
  ram[1350]  = 64;
  ram[1351]  = 0;
  ram[1352]  = 0;
  ram[1353]  = 12;
  ram[1354]  = 226;
  ram[1355]  = 255;
  ram[1356]  = 255;
  ram[1357]  = 255;
  ram[1358]  = 255;
  ram[1359]  = 252;
  ram[1360]  = 244;
  ram[1361]  = 248;
  ram[1362]  = 254;
  ram[1363]  = 253;
  ram[1364]  = 253;
  ram[1365]  = 254;
  ram[1366]  = 253;
  ram[1367]  = 255;
  ram[1368]  = 132;
  ram[1369]  = 0;
  ram[1370]  = 0;
  ram[1371]  = 0;
  ram[1372]  = 0;
  ram[1373]  = 0;
  ram[1374]  = 0;
  ram[1375]  = 1;
  ram[1376]  = 69;
  ram[1377]  = 108;
  ram[1378]  = 137;
  ram[1379]  = 190;
  ram[1380]  = 255;
  ram[1381]  = 183;
  ram[1382]  = 0;
  ram[1383]  = 0;
  ram[1384]  = 0;
  ram[1385]  = 107;
  ram[1386]  = 211;
  ram[1387]  = 10;
  ram[1388]  = 0;
  ram[1389]  = 109;
  ram[1390]  = 255;
  ram[1391]  = 255;
  ram[1392]  = 255;
  ram[1393]  = 255;
  ram[1394]  = 253;
  ram[1395]  = 240;
  ram[1396]  = 252;
  ram[1397]  = 254;
  ram[1398]  = 253;
  ram[1399]  = 254;
  ram[1400]  = 253;
  ram[1401]  = 254;
  ram[1402]  = 253;
  ram[1403]  = 254;
  ram[1404]  = 254;
  ram[1405]  = 250;
  ram[1406]  = 243;
  ram[1407]  = 253;
  ram[1408]  = 255;
  ram[1409]  = 198;
  ram[1410]  = 78;
  ram[1411]  = 38;
  ram[1412]  = 88;
  ram[1413]  = 131;
  ram[1414]  = 127;
  ram[1415]  = 165;
  ram[1416]  = 200;
  ram[1417]  = 218;
  ram[1418]  = 234;
  ram[1419]  = 255;
  ram[1420]  = 164;
  ram[1421]  = 0;
  ram[1422]  = 0;
  ram[1423]  = 0;
  ram[1424]  = 0;
  ram[1425]  = 47;
  ram[1426]  = 249;
  ram[1427]  = 255;
  ram[1428]  = 246;
  ram[1429]  = 246;
  ram[1430]  = 253;
  ram[1431]  = 252;
  ram[1432]  = 252;
  ram[1433]  = 251;
  ram[1434]  = 251;
  ram[1435]  = 250;
  ram[1436]  = 251;
  ram[1437]  = 253;
  ram[1438]  = 254;
  ram[1439]  = 245;
  ram[1440]  = 251;
  ram[1441]  = 252;
  ram[1442]  = 251;
  ram[1443]  = 252;
  ram[1444]  = 252;
  ram[1445]  = 252;
  ram[1446]  = 251;
  ram[1447]  = 252;
  ram[1448]  = 250;
  ram[1449]  = 243;
  ram[1450]  = 252;
  ram[1451]  = 255;
  ram[1452]  = 104;
  ram[1453]  = 0;
  ram[1454]  = 0;
  ram[1455]  = 23;
  ram[1456]  = 202;
  ram[1457]  = 220;
  ram[1458]  = 245;
  ram[1459]  = 255;
  ram[1460]  = 235;
  ram[1461]  = 32;
  ram[1462]  = 0;
  ram[1463]  = 0;
  ram[1464]  = 11;
  ram[1465]  = 216;
  ram[1466]  = 253;
  ram[1467]  = 252;
  ram[1468]  = 255;
  ram[1469]  = 255;
  ram[1470]  = 199;
  ram[1471]  = 5;
  ram[1472]  = 0;
  ram[1473]  = 106;
  ram[1474]  = 238;
  ram[1475]  = 172;
  ram[1476]  = 133;
  ram[1477]  = 180;
  ram[1478]  = 250;
  ram[1479]  = 251;
  ram[1480]  = 238;
  ram[1481]  = 243;
  ram[1482]  = 249;
  ram[1483]  = 247;
  ram[1484]  = 248;
  ram[1485]  = 247;
  ram[1486]  = 255;
  ram[1487]  = 208;
  ram[1488]  = 10;
  ram[1489]  = 0;
  ram[1490]  = 0;
  ram[1491]  = 1;
  ram[1492]  = 128;
  ram[1493]  = 78;
  ram[1494]  = 0;
  ram[1495]  = 1;
  ram[1496]  = 126;
  ram[1497]  = 255;
  ram[1498]  = 255;
  ram[1499]  = 255;
  ram[1500]  = 241;
  ram[1501]  = 52;
  ram[1502]  = 0;
  ram[1503]  = 0;
  ram[1504]  = 7;
  ram[1505]  = 228;
  ram[1506]  = 223;
  ram[1507]  = 0;
  ram[1508]  = 0;
  ram[1509]  = 0;
  ram[1510]  = 66;
  ram[1511]  = 232;
  ram[1512]  = 254;
  ram[1513]  = 249;
  ram[1514]  = 244;
  ram[1515]  = 236;
  ram[1516]  = 245;
  ram[1517]  = 246;
  ram[1518]  = 247;
  ram[1519]  = 248;
  ram[1520]  = 245;
  ram[1521]  = 246;
  ram[1522]  = 248;
  ram[1523]  = 248;
  ram[1524]  = 247;
  ram[1525]  = 242;
  ram[1526]  = 236;
  ram[1527]  = 247;
  ram[1528]  = 247;
  ram[1529]  = 255;
  ram[1530]  = 255;
  ram[1531]  = 239;
  ram[1532]  = 255;
  ram[1533]  = 255;
  ram[1534]  = 255;
  ram[1535]  = 255;
  ram[1536]  = 255;
  ram[1537]  = 247;
  ram[1538]  = 255;
  ram[1539]  = 222;
  ram[1540]  = 22;
  ram[1541]  = 0;
  ram[1542]  = 0;
  ram[1543]  = 0;
  ram[1544]  = 0;
  ram[1545]  = 164;
  ram[1546]  = 255;
  ram[1547]  = 242;
  ram[1548]  = 240;
  ram[1549]  = 238;
  ram[1550]  = 245;
  ram[1551]  = 243;
  ram[1552]  = 242;
  ram[1553]  = 242;
  ram[1554]  = 244;
  ram[1555]  = 242;
  ram[1556]  = 244;
  ram[1557]  = 243;
  ram[1558]  = 244;
  ram[1559]  = 234;
  ram[1560]  = 240;
  ram[1561]  = 239;
  ram[1562]  = 237;
  ram[1563]  = 239;
  ram[1564]  = 237;
  ram[1565]  = 238;
  ram[1566]  = 241;
  ram[1567]  = 244;
  ram[1568]  = 249;
  ram[1569]  = 250;
  ram[1570]  = 255;
  ram[1571]  = 255;
  ram[1572]  = 108;
  ram[1573]  = 0;
  ram[1574]  = 0;
  ram[1575]  = 0;
  ram[1576]  = 5;
  ram[1577]  = 6;
  ram[1578]  = 75;
  ram[1579]  = 253;
  ram[1580]  = 134;
  ram[1581]  = 0;
  ram[1582]  = 0;
  ram[1583]  = 0;
  ram[1584]  = 95;
  ram[1585]  = 255;
  ram[1586]  = 255;
  ram[1587]  = 251;
  ram[1588]  = 224;
  ram[1589]  = 178;
  ram[1590]  = 91;
  ram[1591]  = 3;
  ram[1592]  = 0;
  ram[1593]  = 24;
  ram[1594]  = 21;
  ram[1595]  = 0;
  ram[1596]  = 0;
  ram[1597]  = 0;
  ram[1598]  = 121;
  ram[1599]  = 254;
  ram[1600]  = 232;
  ram[1601]  = 238;
  ram[1602]  = 243;
  ram[1603]  = 242;
  ram[1604]  = 242;
  ram[1605]  = 246;
  ram[1606]  = 247;
  ram[1607]  = 58;
  ram[1608]  = 0;
  ram[1609]  = 0;
  ram[1610]  = 0;
  ram[1611]  = 90;
  ram[1612]  = 255;
  ram[1613]  = 136;
  ram[1614]  = 0;
  ram[1615]  = 0;
  ram[1616]  = 0;
  ram[1617]  = 107;
  ram[1618]  = 252;
  ram[1619]  = 248;
  ram[1620]  = 199;
  ram[1621]  = 0;
  ram[1622]  = 0;
  ram[1623]  = 0;
  ram[1624]  = 100;
  ram[1625]  = 255;
  ram[1626]  = 244;
  ram[1627]  = 82;
  ram[1628]  = 0;
  ram[1629]  = 0;
  ram[1630]  = 0;
  ram[1631]  = 94;
  ram[1632]  = 255;
  ram[1633]  = 242;
  ram[1634]  = 238;
  ram[1635]  = 231;
  ram[1636]  = 240;
  ram[1637]  = 242;
  ram[1638]  = 243;
  ram[1639]  = 243;
  ram[1640]  = 241;
  ram[1641]  = 242;
  ram[1642]  = 242;
  ram[1643]  = 244;
  ram[1644]  = 243;
  ram[1645]  = 237;
  ram[1646]  = 230;
  ram[1647]  = 240;
  ram[1648]  = 241;
  ram[1649]  = 242;
  ram[1650]  = 240;
  ram[1651]  = 243;
  ram[1652]  = 242;
  ram[1653]  = 239;
  ram[1654]  = 241;
  ram[1655]  = 240;
  ram[1656]  = 241;
  ram[1657]  = 236;
  ram[1658]  = 241;
  ram[1659]  = 65;
  ram[1660]  = 0;
  ram[1661]  = 0;
  ram[1662]  = 0;
  ram[1663]  = 0;
  ram[1664]  = 124;
  ram[1665]  = 255;
  ram[1666]  = 246;
  ram[1667]  = 241;
  ram[1668]  = 238;
  ram[1669]  = 237;
  ram[1670]  = 246;
  ram[1671]  = 245;
  ram[1672]  = 244;
  ram[1673]  = 245;
  ram[1674]  = 244;
  ram[1675]  = 242;
  ram[1676]  = 242;
  ram[1677]  = 243;
  ram[1678]  = 245;
  ram[1679]  = 234;
  ram[1680]  = 250;
  ram[1681]  = 247;
  ram[1682]  = 246;
  ram[1683]  = 247;
  ram[1684]  = 247;
  ram[1685]  = 248;
  ram[1686]  = 251;
  ram[1687]  = 255;
  ram[1688]  = 230;
  ram[1689]  = 188;
  ram[1690]  = 112;
  ram[1691]  = 53;
  ram[1692]  = 10;
  ram[1693]  = 0;
  ram[1694]  = 0;
  ram[1695]  = 0;
  ram[1696]  = 0;
  ram[1697]  = 0;
  ram[1698]  = 0;
  ram[1699]  = 181;
  ram[1700]  = 36;
  ram[1701]  = 0;
  ram[1702]  = 0;
  ram[1703]  = 14;
  ram[1704]  = 213;
  ram[1705]  = 214;
  ram[1706]  = 110;
  ram[1707]  = 59;
  ram[1708]  = 22;
  ram[1709]  = 0;
  ram[1710]  = 0;
  ram[1711]  = 0;
  ram[1712]  = 0;
  ram[1713]  = 0;
  ram[1714]  = 0;
  ram[1715]  = 0;
  ram[1716]  = 0;
  ram[1717]  = 0;
  ram[1718]  = 67;
  ram[1719]  = 253;
  ram[1720]  = 243;
  ram[1721]  = 247;
  ram[1722]  = 253;
  ram[1723]  = 252;
  ram[1724]  = 252;
  ram[1725]  = 255;
  ram[1726]  = 167;
  ram[1727]  = 0;
  ram[1728]  = 0;
  ram[1729]  = 0;
  ram[1730]  = 32;
  ram[1731]  = 229;
  ram[1732]  = 251;
  ram[1733]  = 229;
  ram[1734]  = 51;
  ram[1735]  = 0;
  ram[1736]  = 0;
  ram[1737]  = 0;
  ram[1738]  = 170;
  ram[1739]  = 255;
  ram[1740]  = 232;
  ram[1741]  = 40;
  ram[1742]  = 0;
  ram[1743]  = 46;
  ram[1744]  = 236;
  ram[1745]  = 254;
  ram[1746]  = 255;
  ram[1747]  = 252;
  ram[1748]  = 90;
  ram[1749]  = 0;
  ram[1750]  = 0;
  ram[1751]  = 122;
  ram[1752]  = 255;
  ram[1753]  = 252;
  ram[1754]  = 247;
  ram[1755]  = 241;
  ram[1756]  = 251;
  ram[1757]  = 252;
  ram[1758]  = 253;
  ram[1759]  = 252;
  ram[1760]  = 251;
  ram[1761]  = 252;
  ram[1762]  = 253;
  ram[1763]  = 253;
  ram[1764]  = 254;
  ram[1765]  = 246;
  ram[1766]  = 240;
  ram[1767]  = 250;
  ram[1768]  = 251;
  ram[1769]  = 251;
  ram[1770]  = 252;
  ram[1771]  = 251;
  ram[1772]  = 251;
  ram[1773]  = 249;
  ram[1774]  = 251;
  ram[1775]  = 252;
  ram[1776]  = 255;
  ram[1777]  = 255;
  ram[1778]  = 119;
  ram[1779]  = 0;
  ram[1780]  = 0;
  ram[1781]  = 0;
  ram[1782]  = 0;
  ram[1783]  = 82;
  ram[1784]  = 254;
  ram[1785]  = 254;
  ram[1786]  = 252;
  ram[1787]  = 251;
  ram[1788]  = 245;
  ram[1789]  = 245;
  ram[1790]  = 253;
  ram[1791]  = 253;
  ram[1792]  = 252;
  ram[1793]  = 252;
  ram[1794]  = 250;
  ram[1795]  = 251;
  ram[1796]  = 251;
  ram[1797]  = 252;
  ram[1798]  = 254;
  ram[1799]  = 244;
  ram[1800]  = 252;
  ram[1801]  = 251;
  ram[1802]  = 253;
  ram[1803]  = 253;
  ram[1804]  = 251;
  ram[1805]  = 253;
  ram[1806]  = 255;
  ram[1807]  = 146;
  ram[1808]  = 24;
  ram[1809]  = 0;
  ram[1810]  = 0;
  ram[1811]  = 0;
  ram[1812]  = 0;
  ram[1813]  = 0;
  ram[1814]  = 0;
  ram[1815]  = 0;
  ram[1816]  = 0;
  ram[1817]  = 0;
  ram[1818]  = 79;
  ram[1819]  = 116;
  ram[1820]  = 0;
  ram[1821]  = 0;
  ram[1822]  = 0;
  ram[1823]  = 37;
  ram[1824]  = 247;
  ram[1825]  = 51;
  ram[1826]  = 0;
  ram[1827]  = 0;
  ram[1828]  = 0;
  ram[1829]  = 0;
  ram[1830]  = 0;
  ram[1831]  = 0;
  ram[1832]  = 0;
  ram[1833]  = 0;
  ram[1834]  = 0;
  ram[1835]  = 3;
  ram[1836]  = 20;
  ram[1837]  = 74;
  ram[1838]  = 232;
  ram[1839]  = 254;
  ram[1840]  = 241;
  ram[1841]  = 247;
  ram[1842]  = 253;
  ram[1843]  = 252;
  ram[1844]  = 252;
  ram[1845]  = 255;
  ram[1846]  = 121;
  ram[1847]  = 0;
  ram[1848]  = 0;
  ram[1849]  = 13;
  ram[1850]  = 200;
  ram[1851]  = 255;
  ram[1852]  = 242;
  ram[1853]  = 255;
  ram[1854]  = 229;
  ram[1855]  = 41;
  ram[1856]  = 0;
  ram[1857]  = 0;
  ram[1858]  = 141;
  ram[1859]  = 255;
  ram[1860]  = 255;
  ram[1861]  = 221;
  ram[1862]  = 171;
  ram[1863]  = 220;
  ram[1864]  = 255;
  ram[1865]  = 252;
  ram[1866]  = 252;
  ram[1867]  = 255;
  ram[1868]  = 255;
  ram[1869]  = 169;
  ram[1870]  = 157;
  ram[1871]  = 255;
  ram[1872]  = 255;
  ram[1873]  = 252;
  ram[1874]  = 247;
  ram[1875]  = 242;
  ram[1876]  = 253;
  ram[1877]  = 253;
  ram[1878]  = 252;
  ram[1879]  = 252;
  ram[1880]  = 252;
  ram[1881]  = 252;
  ram[1882]  = 253;
  ram[1883]  = 252;
  ram[1884]  = 253;
  ram[1885]  = 247;
  ram[1886]  = 240;
  ram[1887]  = 251;
  ram[1888]  = 251;
  ram[1889]  = 252;
  ram[1890]  = 251;
  ram[1891]  = 251;
  ram[1892]  = 251;
  ram[1893]  = 250;
  ram[1894]  = 252;
  ram[1895]  = 254;
  ram[1896]  = 255;
  ram[1897]  = 153;
  ram[1898]  = 0;
  ram[1899]  = 0;
  ram[1900]  = 0;
  ram[1901]  = 0;
  ram[1902]  = 53;
  ram[1903]  = 239;
  ram[1904]  = 255;
  ram[1905]  = 252;
  ram[1906]  = 252;
  ram[1907]  = 252;
  ram[1908]  = 246;
  ram[1909]  = 242;
  ram[1910]  = 253;
  ram[1911]  = 252;
  ram[1912]  = 252;
  ram[1913]  = 252;
  ram[1914]  = 250;
  ram[1915]  = 252;
  ram[1916]  = 252;
  ram[1917]  = 251;
  ram[1918]  = 253;
  ram[1919]  = 244;
  ram[1920]  = 250;
  ram[1921]  = 249;
  ram[1922]  = 251;
  ram[1923]  = 252;
  ram[1924]  = 252;
  ram[1925]  = 253;
  ram[1926]  = 255;
  ram[1927]  = 58;
  ram[1928]  = 0;
  ram[1929]  = 0;
  ram[1930]  = 0;
  ram[1931]  = 0;
  ram[1932]  = 0;
  ram[1933]  = 0;
  ram[1934]  = 0;
  ram[1935]  = 0;
  ram[1936]  = 50;
  ram[1937]  = 130;
  ram[1938]  = 227;
  ram[1939]  = 29;
  ram[1940]  = 0;
  ram[1941]  = 0;
  ram[1942]  = 0;
  ram[1943]  = 0;
  ram[1944]  = 207;
  ram[1945]  = 120;
  ram[1946]  = 0;
  ram[1947]  = 0;
  ram[1948]  = 0;
  ram[1949]  = 15;
  ram[1950]  = 4;
  ram[1951]  = 0;
  ram[1952]  = 0;
  ram[1953]  = 78;
  ram[1954]  = 181;
  ram[1955]  = 210;
  ram[1956]  = 231;
  ram[1957]  = 255;
  ram[1958]  = 255;
  ram[1959]  = 252;
  ram[1960]  = 244;
  ram[1961]  = 248;
  ram[1962]  = 251;
  ram[1963]  = 252;
  ram[1964]  = 252;
  ram[1965]  = 254;
  ram[1966]  = 201;
  ram[1967]  = 70;
  ram[1968]  = 35;
  ram[1969]  = 178;
  ram[1970]  = 255;
  ram[1971]  = 249;
  ram[1972]  = 247;
  ram[1973]  = 255;
  ram[1974]  = 255;
  ram[1975]  = 228;
  ram[1976]  = 77;
  ram[1977]  = 122;
  ram[1978]  = 230;
  ram[1979]  = 254;
  ram[1980]  = 251;
  ram[1981]  = 255;
  ram[1982]  = 255;
  ram[1983]  = 246;
  ram[1984]  = 255;
  ram[1985]  = 255;
  ram[1986]  = 255;
  ram[1987]  = 248;
  ram[1988]  = 217;
  ram[1989]  = 209;
  ram[1990]  = 237;
  ram[1991]  = 234;
  ram[1992]  = 255;
  ram[1993]  = 255;
  ram[1994]  = 246;
  ram[1995]  = 242;
  ram[1996]  = 253;
  ram[1997]  = 251;
  ram[1998]  = 251;
  ram[1999]  = 252;
  ram[2000]  = 253;
  ram[2001]  = 253;
  ram[2002]  = 252;
  ram[2003]  = 251;
  ram[2004]  = 252;
  ram[2005]  = 248;
  ram[2006]  = 240;
  ram[2007]  = 252;
  ram[2008]  = 253;
  ram[2009]  = 252;
  ram[2010]  = 251;
  ram[2011]  = 252;
  ram[2012]  = 252;
  ram[2013]  = 252;
  ram[2014]  = 252;
  ram[2015]  = 255;
  ram[2016]  = 184;
  ram[2017]  = 5;
  ram[2018]  = 0;
  ram[2019]  = 0;
  ram[2020]  = 0;
  ram[2021]  = 27;
  ram[2022]  = 222;
  ram[2023]  = 255;
  ram[2024]  = 252;
  ram[2025]  = 252;
  ram[2026]  = 252;
  ram[2027]  = 253;
  ram[2028]  = 247;
  ram[2029]  = 244;
  ram[2030]  = 253;
  ram[2031]  = 252;
  ram[2032]  = 253;
  ram[2033]  = 252;
  ram[2034]  = 251;
  ram[2035]  = 252;
  ram[2036]  = 252;
  ram[2037]  = 253;
  ram[2038]  = 253;
  ram[2039]  = 245;
  ram[2040]  = 252;
  ram[2041]  = 251;
  ram[2042]  = 250;
  ram[2043]  = 250;
  ram[2044]  = 251;
  ram[2045]  = 252;
  ram[2046]  = 255;
  ram[2047]  = 205;
  ram[2048]  = 53;
  ram[2049]  = 0;
  ram[2050]  = 7;
  ram[2051]  = 40;
  ram[2052]  = 33;
  ram[2053]  = 0;
  ram[2054]  = 0;
  ram[2055]  = 0;
  ram[2056]  = 196;
  ram[2057]  = 255;
  ram[2058]  = 116;
  ram[2059]  = 0;
  ram[2060]  = 0;
  ram[2061]  = 0;
  ram[2062]  = 0;
  ram[2063]  = 0;
  ram[2064]  = 178;
  ram[2065]  = 253;
  ram[2066]  = 181;
  ram[2067]  = 151;
  ram[2068]  = 197;
  ram[2069]  = 219;
  ram[2070]  = 32;
  ram[2071]  = 0;
  ram[2072]  = 0;
  ram[2073]  = 152;
  ram[2074]  = 255;
  ram[2075]  = 255;
  ram[2076]  = 255;
  ram[2077]  = 253;
  ram[2078]  = 252;
  ram[2079]  = 252;
  ram[2080]  = 244;
  ram[2081]  = 248;
  ram[2082]  = 252;
  ram[2083]  = 253;
  ram[2084]  = 252;
  ram[2085]  = 251;
  ram[2086]  = 255;
  ram[2087]  = 255;
  ram[2088]  = 245;
  ram[2089]  = 255;
  ram[2090]  = 254;
  ram[2091]  = 251;
  ram[2092]  = 246;
  ram[2093]  = 107;
  ram[2094]  = 61;
  ram[2095]  = 192;
  ram[2096]  = 255;
  ram[2097]  = 255;
  ram[2098]  = 255;
  ram[2099]  = 252;
  ram[2100]  = 251;
  ram[2101]  = 253;
  ram[2102]  = 255;
  ram[2103]  = 255;
  ram[2104]  = 231;
  ram[2105]  = 173;
  ram[2106]  = 106;
  ram[2107]  = 43;
  ram[2108]  = 7;
  ram[2109]  = 0;
  ram[2110]  = 11;
  ram[2111]  = 20;
  ram[2112]  = 99;
  ram[2113]  = 239;
  ram[2114]  = 255;
  ram[2115]  = 242;
  ram[2116]  = 252;
  ram[2117]  = 252;
  ram[2118]  = 252;
  ram[2119]  = 252;
  ram[2120]  = 252;
  ram[2121]  = 253;
  ram[2122]  = 252;
  ram[2123]  = 252;
  ram[2124]  = 253;
  ram[2125]  = 248;
  ram[2126]  = 242;
  ram[2127]  = 253;
  ram[2128]  = 252;
  ram[2129]  = 252;
  ram[2130]  = 253;
  ram[2131]  = 252;
  ram[2132]  = 252;
  ram[2133]  = 252;
  ram[2134]  = 255;
  ram[2135]  = 237;
  ram[2136]  = 29;
  ram[2137]  = 0;
  ram[2138]  = 0;
  ram[2139]  = 0;
  ram[2140]  = 30;
  ram[2141]  = 201;
  ram[2142]  = 255;
  ram[2143]  = 253;
  ram[2144]  = 253;
  ram[2145]  = 253;
  ram[2146]  = 253;
  ram[2147]  = 253;
  ram[2148]  = 250;
  ram[2149]  = 250;
  ram[2150]  = 253;
  ram[2151]  = 255;
  ram[2152]  = 255;
  ram[2153]  = 253;
  ram[2154]  = 252;
  ram[2155]  = 252;
  ram[2156]  = 252;
  ram[2157]  = 251;
  ram[2158]  = 253;
  ram[2159]  = 246;
  ram[2160]  = 250;
  ram[2161]  = 252;
  ram[2162]  = 252;
  ram[2163]  = 249;
  ram[2164]  = 249;
  ram[2165]  = 251;
  ram[2166]  = 251;
  ram[2167]  = 255;
  ram[2168]  = 248;
  ram[2169]  = 196;
  ram[2170]  = 215;
  ram[2171]  = 249;
  ram[2172]  = 174;
  ram[2173]  = 0;
  ram[2174]  = 0;
  ram[2175]  = 0;
  ram[2176]  = 201;
  ram[2177]  = 235;
  ram[2178]  = 7;
  ram[2179]  = 0;
  ram[2180]  = 0;
  ram[2181]  = 0;
  ram[2182]  = 0;
  ram[2183]  = 0;
  ram[2184]  = 176;
  ram[2185]  = 255;
  ram[2186]  = 255;
  ram[2187]  = 255;
  ram[2188]  = 255;
  ram[2189]  = 248;
  ram[2190]  = 28;
  ram[2191]  = 0;
  ram[2192]  = 0;
  ram[2193]  = 116;
  ram[2194]  = 255;
  ram[2195]  = 251;
  ram[2196]  = 255;
  ram[2197]  = 255;
  ram[2198]  = 251;
  ram[2199]  = 251;
  ram[2200]  = 245;
  ram[2201]  = 250;
  ram[2202]  = 252;
  ram[2203]  = 252;
  ram[2204]  = 252;
  ram[2205]  = 252;
  ram[2206]  = 252;
  ram[2207]  = 255;
  ram[2208]  = 255;
  ram[2209]  = 254;
  ram[2210]  = 254;
  ram[2211]  = 255;
  ram[2212]  = 220;
  ram[2213]  = 6;
  ram[2214]  = 0;
  ram[2215]  = 75;
  ram[2216]  = 255;
  ram[2217]  = 254;
  ram[2218]  = 253;
  ram[2219]  = 253;
  ram[2220]  = 252;
  ram[2221]  = 254;
  ram[2222]  = 197;
  ram[2223]  = 127;
  ram[2224]  = 24;
  ram[2225]  = 0;
  ram[2226]  = 0;
  ram[2227]  = 0;
  ram[2228]  = 0;
  ram[2229]  = 0;
  ram[2230]  = 0;
  ram[2231]  = 0;
  ram[2232]  = 0;
  ram[2233]  = 47;
  ram[2234]  = 235;
  ram[2235]  = 251;
  ram[2236]  = 253;
  ram[2237]  = 252;
  ram[2238]  = 250;
  ram[2239]  = 252;
  ram[2240]  = 252;
  ram[2241]  = 252;
  ram[2242]  = 252;
  ram[2243]  = 253;
  ram[2244]  = 253;
  ram[2245]  = 248;
  ram[2246]  = 244;
  ram[2247]  = 253;
  ram[2248]  = 252;
  ram[2249]  = 252;
  ram[2250]  = 252;
  ram[2251]  = 252;
  ram[2252]  = 253;
  ram[2253]  = 252;
  ram[2254]  = 255;
  ram[2255]  = 234;
  ram[2256]  = 21;
  ram[2257]  = 0;
  ram[2258]  = 0;
  ram[2259]  = 0;
  ram[2260]  = 108;
  ram[2261]  = 255;
  ram[2262]  = 255;
  ram[2263]  = 255;
  ram[2264]  = 255;
  ram[2265]  = 255;
  ram[2266]  = 255;
  ram[2267]  = 255;
  ram[2268]  = 255;
  ram[2269]  = 255;
  ram[2270]  = 255;
  ram[2271]  = 255;
  ram[2272]  = 255;
  ram[2273]  = 255;
  ram[2274]  = 254;
  ram[2275]  = 253;
  ram[2276]  = 252;
  ram[2277]  = 251;
  ram[2278]  = 252;
  ram[2279]  = 244;
  ram[2280]  = 250;
  ram[2281]  = 250;
  ram[2282]  = 252;
  ram[2283]  = 250;
  ram[2284]  = 251;
  ram[2285]  = 251;
  ram[2286]  = 249;
  ram[2287]  = 249;
  ram[2288]  = 252;
  ram[2289]  = 255;
  ram[2290]  = 255;
  ram[2291]  = 255;
  ram[2292]  = 177;
  ram[2293]  = 0;
  ram[2294]  = 0;
  ram[2295]  = 0;
  ram[2296]  = 200;
  ram[2297]  = 243;
  ram[2298]  = 14;
  ram[2299]  = 0;
  ram[2300]  = 4;
  ram[2301]  = 15;
  ram[2302]  = 0;
  ram[2303]  = 0;
  ram[2304]  = 180;
  ram[2305]  = 255;
  ram[2306]  = 255;
  ram[2307]  = 255;
  ram[2308]  = 255;
  ram[2309]  = 240;
  ram[2310]  = 34;
  ram[2311]  = 0;
  ram[2312]  = 0;
  ram[2313]  = 45;
  ram[2314]  = 92;
  ram[2315]  = 45;
  ram[2316]  = 81;
  ram[2317]  = 219;
  ram[2318]  = 255;
  ram[2319]  = 251;
  ram[2320]  = 246;
  ram[2321]  = 250;
  ram[2322]  = 252;
  ram[2323]  = 251;
  ram[2324]  = 252;
  ram[2325]  = 250;
  ram[2326]  = 251;
  ram[2327]  = 253;
  ram[2328]  = 253;
  ram[2329]  = 253;
  ram[2330]  = 254;
  ram[2331]  = 255;
  ram[2332]  = 210;
  ram[2333]  = 14;
  ram[2334]  = 0;
  ram[2335]  = 45;
  ram[2336]  = 255;
  ram[2337]  = 255;
  ram[2338]  = 255;
  ram[2339]  = 255;
  ram[2340]  = 255;
  ram[2341]  = 180;
  ram[2342]  = 0;
  ram[2343]  = 0;
  ram[2344]  = 0;
  ram[2345]  = 0;
  ram[2346]  = 0;
  ram[2347]  = 0;
  ram[2348]  = 0;
  ram[2349]  = 19;
  ram[2350]  = 5;
  ram[2351]  = 0;
  ram[2352]  = 0;
  ram[2353]  = 0;
  ram[2354]  = 164;
  ram[2355]  = 255;
  ram[2356]  = 253;
  ram[2357]  = 253;
  ram[2358]  = 251;
  ram[2359]  = 252;
  ram[2360]  = 252;
  ram[2361]  = 252;
  ram[2362]  = 251;
  ram[2363]  = 253;
  ram[2364]  = 253;
  ram[2365]  = 248;
  ram[2366]  = 243;
  ram[2367]  = 252;
  ram[2368]  = 251;
  ram[2369]  = 253;
  ram[2370]  = 252;
  ram[2371]  = 253;
  ram[2372]  = 254;
  ram[2373]  = 255;
  ram[2374]  = 255;
  ram[2375]  = 255;
  ram[2376]  = 171;
  ram[2377]  = 1;
  ram[2378]  = 0;
  ram[2379]  = 0;
  ram[2380]  = 14;
  ram[2381]  = 203;
  ram[2382]  = 255;
  ram[2383]  = 249;
  ram[2384]  = 230;
  ram[2385]  = 199;
  ram[2386]  = 194;
  ram[2387]  = 171;
  ram[2388]  = 136;
  ram[2389]  = 123;
  ram[2390]  = 110;
  ram[2391]  = 58;
  ram[2392]  = 91;
  ram[2393]  = 207;
  ram[2394]  = 255;
  ram[2395]  = 254;
  ram[2396]  = 252;
  ram[2397]  = 251;
  ram[2398]  = 251;
  ram[2399]  = 246;
  ram[2400]  = 251;
  ram[2401]  = 250;
  ram[2402]  = 251;
  ram[2403]  = 251;
  ram[2404]  = 251;
  ram[2405]  = 251;
  ram[2406]  = 249;
  ram[2407]  = 249;
  ram[2408]  = 248;
  ram[2409]  = 241;
  ram[2410]  = 252;
  ram[2411]  = 255;
  ram[2412]  = 169;
  ram[2413]  = 0;
  ram[2414]  = 0;
  ram[2415]  = 0;
  ram[2416]  = 143;
  ram[2417]  = 208;
  ram[2418]  = 180;
  ram[2419]  = 87;
  ram[2420]  = 158;
  ram[2421]  = 56;
  ram[2422]  = 0;
  ram[2423]  = 0;
  ram[2424]  = 152;
  ram[2425]  = 255;
  ram[2426]  = 181;
  ram[2427]  = 131;
  ram[2428]  = 94;
  ram[2429]  = 37;
  ram[2430]  = 2;
  ram[2431]  = 0;
  ram[2432]  = 0;
  ram[2433]  = 0;
  ram[2434]  = 0;
  ram[2435]  = 0;
  ram[2436]  = 0;
  ram[2437]  = 38;
  ram[2438]  = 239;
  ram[2439]  = 254;
  ram[2440]  = 241;
  ram[2441]  = 248;
  ram[2442]  = 252;
  ram[2443]  = 251;
  ram[2444]  = 251;
  ram[2445]  = 250;
  ram[2446]  = 252;
  ram[2447]  = 253;
  ram[2448]  = 253;
  ram[2449]  = 255;
  ram[2450]  = 255;
  ram[2451]  = 255;
  ram[2452]  = 213;
  ram[2453]  = 3;
  ram[2454]  = 0;
  ram[2455]  = 23;
  ram[2456]  = 130;
  ram[2457]  = 125;
  ram[2458]  = 179;
  ram[2459]  = 248;
  ram[2460]  = 255;
  ram[2461]  = 119;
  ram[2462]  = 0;
  ram[2463]  = 1;
  ram[2464]  = 71;
  ram[2465]  = 89;
  ram[2466]  = 129;
  ram[2467]  = 170;
  ram[2468]  = 197;
  ram[2469]  = 234;
  ram[2470]  = 201;
  ram[2471]  = 17;
  ram[2472]  = 0;
  ram[2473]  = 0;
  ram[2474]  = 89;
  ram[2475]  = 255;
  ram[2476]  = 252;
  ram[2477]  = 254;
  ram[2478]  = 253;
  ram[2479]  = 252;
  ram[2480]  = 252;
  ram[2481]  = 252;
  ram[2482]  = 252;
  ram[2483]  = 252;
  ram[2484]  = 253;
  ram[2485]  = 249;
  ram[2486]  = 246;
  ram[2487]  = 255;
  ram[2488]  = 255;
  ram[2489]  = 255;
  ram[2490]  = 255;
  ram[2491]  = 255;
  ram[2492]  = 255;
  ram[2493]  = 246;
  ram[2494]  = 239;
  ram[2495]  = 223;
  ram[2496]  = 165;
  ram[2497]  = 6;
  ram[2498]  = 0;
  ram[2499]  = 0;
  ram[2500]  = 0;
  ram[2501]  = 20;
  ram[2502]  = 58;
  ram[2503]  = 43;
  ram[2504]  = 22;
  ram[2505]  = 0;
  ram[2506]  = 0;
  ram[2507]  = 0;
  ram[2508]  = 0;
  ram[2509]  = 0;
  ram[2510]  = 0;
  ram[2511]  = 0;
  ram[2512]  = 0;
  ram[2513]  = 2;
  ram[2514]  = 168;
  ram[2515]  = 255;
  ram[2516]  = 252;
  ram[2517]  = 251;
  ram[2518]  = 252;
  ram[2519]  = 246;
  ram[2520]  = 252;
  ram[2521]  = 252;
  ram[2522]  = 253;
  ram[2523]  = 250;
  ram[2524]  = 250;
  ram[2525]  = 250;
  ram[2526]  = 250;
  ram[2527]  = 250;
  ram[2528]  = 247;
  ram[2529]  = 241;
  ram[2530]  = 251;
  ram[2531]  = 255;
  ram[2532]  = 199;
  ram[2533]  = 1;
  ram[2534]  = 0;
  ram[2535]  = 1;
  ram[2536]  = 17;
  ram[2537]  = 0;
  ram[2538]  = 95;
  ram[2539]  = 255;
  ram[2540]  = 255;
  ram[2541]  = 55;
  ram[2542]  = 0;
  ram[2543]  = 0;
  ram[2544]  = 177;
  ram[2545]  = 210;
  ram[2546]  = 0;
  ram[2547]  = 0;
  ram[2548]  = 0;
  ram[2549]  = 0;
  ram[2550]  = 0;
  ram[2551]  = 0;
  ram[2552]  = 0;
  ram[2553]  = 0;
  ram[2554]  = 0;
  ram[2555]  = 0;
  ram[2556]  = 0;
  ram[2557]  = 96;
  ram[2558]  = 250;
  ram[2559]  = 252;
  ram[2560]  = 239;
  ram[2561]  = 246;
  ram[2562]  = 253;
  ram[2563]  = 251;
  ram[2564]  = 250;
  ram[2565]  = 251;
  ram[2566]  = 254;
  ram[2567]  = 255;
  ram[2568]  = 255;
  ram[2569]  = 255;
  ram[2570]  = 219;
  ram[2571]  = 173;
  ram[2572]  = 80;
  ram[2573]  = 0;
  ram[2574]  = 0;
  ram[2575]  = 0;
  ram[2576]  = 0;
  ram[2577]  = 0;
  ram[2578]  = 0;
  ram[2579]  = 131;
  ram[2580]  = 255;
  ram[2581]  = 101;
  ram[2582]  = 0;
  ram[2583]  = 0;
  ram[2584]  = 98;
  ram[2585]  = 255;
  ram[2586]  = 255;
  ram[2587]  = 255;
  ram[2588]  = 255;
  ram[2589]  = 255;
  ram[2590]  = 255;
  ram[2591]  = 53;
  ram[2592]  = 0;
  ram[2593]  = 0;
  ram[2594]  = 53;
  ram[2595]  = 253;
  ram[2596]  = 255;
  ram[2597]  = 253;
  ram[2598]  = 253;
  ram[2599]  = 253;
  ram[2600]  = 252;
  ram[2601]  = 252;
  ram[2602]  = 254;
  ram[2603]  = 255;
  ram[2604]  = 255;
  ram[2605]  = 255;
  ram[2606]  = 255;
  ram[2607]  = 254;
  ram[2608]  = 234;
  ram[2609]  = 207;
  ram[2610]  = 162;
  ram[2611]  = 113;
  ram[2612]  = 84;
  ram[2613]  = 39;
  ram[2614]  = 27;
  ram[2615]  = 12;
  ram[2616]  = 0;
  ram[2617]  = 0;
  ram[2618]  = 0;
  ram[2619]  = 0;
  ram[2620]  = 0;
  ram[2621]  = 0;
  ram[2622]  = 0;
  ram[2623]  = 0;
  ram[2624]  = 0;
  ram[2625]  = 0;
  ram[2626]  = 0;
  ram[2627]  = 0;
  ram[2628]  = 0;
  ram[2629]  = 0;
  ram[2630]  = 0;
  ram[2631]  = 0;
  ram[2632]  = 0;
  ram[2633]  = 0;
  ram[2634]  = 52;
  ram[2635]  = 247;
  ram[2636]  = 252;
  ram[2637]  = 251;
  ram[2638]  = 252;
  ram[2639]  = 248;
  ram[2640]  = 253;
  ram[2641]  = 252;
  ram[2642]  = 251;
  ram[2643]  = 252;
  ram[2644]  = 251;
  ram[2645]  = 251;
  ram[2646]  = 251;
  ram[2647]  = 252;
  ram[2648]  = 249;
  ram[2649]  = 243;
  ram[2650]  = 255;
  ram[2651]  = 255;
  ram[2652]  = 193;
  ram[2653]  = 1;
  ram[2654]  = 0;
  ram[2655]  = 0;
  ram[2656]  = 0;
  ram[2657]  = 0;
  ram[2658]  = 76;
  ram[2659]  = 255;
  ram[2660]  = 245;
  ram[2661]  = 37;
  ram[2662]  = 0;
  ram[2663]  = 0;
  ram[2664]  = 173;
  ram[2665]  = 223;
  ram[2666]  = 29;
  ram[2667]  = 0;
  ram[2668]  = 0;
  ram[2669]  = 0;
  ram[2670]  = 0;
  ram[2671]  = 0;
  ram[2672]  = 0;
  ram[2673]  = 27;
  ram[2674]  = 106;
  ram[2675]  = 134;
  ram[2676]  = 174;
  ram[2677]  = 255;
  ram[2678]  = 253;
  ram[2679]  = 250;
  ram[2680]  = 238;
  ram[2681]  = 248;
  ram[2682]  = 252;
  ram[2683]  = 252;
  ram[2684]  = 252;
  ram[2685]  = 252;
  ram[2686]  = 255;
  ram[2687]  = 200;
  ram[2688]  = 115;
  ram[2689]  = 48;
  ram[2690]  = 9;
  ram[2691]  = 0;
  ram[2692]  = 0;
  ram[2693]  = 0;
  ram[2694]  = 0;
  ram[2695]  = 0;
  ram[2696]  = 0;
  ram[2697]  = 0;
  ram[2698]  = 0;
  ram[2699]  = 134;
  ram[2700]  = 255;
  ram[2701]  = 107;
  ram[2702]  = 0;
  ram[2703]  = 0;
  ram[2704]  = 63;
  ram[2705]  = 255;
  ram[2706]  = 255;
  ram[2707]  = 255;
  ram[2708]  = 255;
  ram[2709]  = 255;
  ram[2710]  = 251;
  ram[2711]  = 68;
  ram[2712]  = 0;
  ram[2713]  = 0;
  ram[2714]  = 24;
  ram[2715]  = 233;
  ram[2716]  = 255;
  ram[2717]  = 253;
  ram[2718]  = 253;
  ram[2719]  = 254;
  ram[2720]  = 253;
  ram[2721]  = 253;
  ram[2722]  = 255;
  ram[2723]  = 236;
  ram[2724]  = 174;
  ram[2725]  = 109;
  ram[2726]  = 83;
  ram[2727]  = 48;
  ram[2728]  = 18;
  ram[2729]  = 3;
  ram[2730]  = 0;
  ram[2731]  = 0;
  ram[2732]  = 0;
  ram[2733]  = 0;
  ram[2734]  = 0;
  ram[2735]  = 0;
  ram[2736]  = 0;
  ram[2737]  = 0;
  ram[2738]  = 0;
  ram[2739]  = 0;
  ram[2740]  = 0;
  ram[2741]  = 0;
  ram[2742]  = 0;
  ram[2743]  = 0;
  ram[2744]  = 0;
  ram[2745]  = 0;
  ram[2746]  = 0;
  ram[2747]  = 0;
  ram[2748]  = 0;
  ram[2749]  = 0;
  ram[2750]  = 0;
  ram[2751]  = 0;
  ram[2752]  = 0;
  ram[2753]  = 0;
  ram[2754]  = 152;
  ram[2755]  = 250;
  ram[2756]  = 254;
  ram[2757]  = 252;
  ram[2758]  = 253;
  ram[2759]  = 246;
  ram[2760]  = 253;
  ram[2761]  = 252;
  ram[2762]  = 252;
  ram[2763]  = 252;
  ram[2764]  = 253;
  ram[2765]  = 253;
  ram[2766]  = 252;
  ram[2767]  = 252;
  ram[2768]  = 253;
  ram[2769]  = 255;
  ram[2770]  = 255;
  ram[2771]  = 158;
  ram[2772]  = 32;
  ram[2773]  = 0;
  ram[2774]  = 0;
  ram[2775]  = 0;
  ram[2776]  = 0;
  ram[2777]  = 0;
  ram[2778]  = 191;
  ram[2779]  = 255;
  ram[2780]  = 236;
  ram[2781]  = 25;
  ram[2782]  = 0;
  ram[2783]  = 0;
  ram[2784]  = 154;
  ram[2785]  = 255;
  ram[2786]  = 233;
  ram[2787]  = 126;
  ram[2788]  = 130;
  ram[2789]  = 160;
  ram[2790]  = 22;
  ram[2791]  = 0;
  ram[2792]  = 0;
  ram[2793]  = 93;
  ram[2794]  = 255;
  ram[2795]  = 255;
  ram[2796]  = 255;
  ram[2797]  = 253;
  ram[2798]  = 252;
  ram[2799]  = 251;
  ram[2800]  = 236;
  ram[2801]  = 248;
  ram[2802]  = 254;
  ram[2803]  = 252;
  ram[2804]  = 252;
  ram[2805]  = 255;
  ram[2806]  = 191;
  ram[2807]  = 0;
  ram[2808]  = 0;
  ram[2809]  = 0;
  ram[2810]  = 0;
  ram[2811]  = 0;
  ram[2812]  = 0;
  ram[2813]  = 0;
  ram[2814]  = 0;
  ram[2815]  = 0;
  ram[2816]  = 0;
  ram[2817]  = 29;
  ram[2818]  = 138;
  ram[2819]  = 244;
  ram[2820]  = 255;
  ram[2821]  = 95;
  ram[2822]  = 0;
  ram[2823]  = 0;
  ram[2824]  = 42;
  ram[2825]  = 199;
  ram[2826]  = 152;
  ram[2827]  = 106;
  ram[2828]  = 70;
  ram[2829]  = 62;
  ram[2830]  = 39;
  ram[2831]  = 10;
  ram[2832]  = 0;
  ram[2833]  = 0;
  ram[2834]  = 6;
  ram[2835]  = 215;
  ram[2836]  = 255;
  ram[2837]  = 253;
  ram[2838]  = 253;
  ram[2839]  = 253;
  ram[2840]  = 254;
  ram[2841]  = 255;
  ram[2842]  = 158;
  ram[2843]  = 33;
  ram[2844]  = 0;
  ram[2845]  = 0;
  ram[2846]  = 0;
  ram[2847]  = 0;
  ram[2848]  = 0;
  ram[2849]  = 0;
  ram[2850]  = 0;
  ram[2851]  = 0;
  ram[2852]  = 0;
  ram[2853]  = 0;
  ram[2854]  = 0;
  ram[2855]  = 0;
  ram[2856]  = 0;
  ram[2857]  = 0;
  ram[2858]  = 0;
  ram[2859]  = 0;
  ram[2860]  = 0;
  ram[2861]  = 0;
  ram[2862]  = 0;
  ram[2863]  = 0;
  ram[2864]  = 11;
  ram[2865]  = 32;
  ram[2866]  = 56;
  ram[2867]  = 96;
  ram[2868]  = 81;
  ram[2869]  = 74;
  ram[2870]  = 80;
  ram[2871]  = 100;
  ram[2872]  = 87;
  ram[2873]  = 170;
  ram[2874]  = 255;
  ram[2875]  = 255;
  ram[2876]  = 252;
  ram[2877]  = 253;
  ram[2878]  = 253;
  ram[2879]  = 248;
  ram[2880]  = 253;
  ram[2881]  = 253;
  ram[2882]  = 253;
  ram[2883]  = 253;
  ram[2884]  = 254;
  ram[2885]  = 253;
  ram[2886]  = 253;
  ram[2887]  = 255;
  ram[2888]  = 255;
  ram[2889]  = 196;
  ram[2890]  = 65;
  ram[2891]  = 0;
  ram[2892]  = 0;
  ram[2893]  = 0;
  ram[2894]  = 0;
  ram[2895]  = 0;
  ram[2896]  = 18;
  ram[2897]  = 170;
  ram[2898]  = 255;
  ram[2899]  = 255;
  ram[2900]  = 224;
  ram[2901]  = 13;
  ram[2902]  = 0;
  ram[2903]  = 0;
  ram[2904]  = 159;
  ram[2905]  = 255;
  ram[2906]  = 255;
  ram[2907]  = 255;
  ram[2908]  = 255;
  ram[2909]  = 255;
  ram[2910]  = 32;
  ram[2911]  = 0;
  ram[2912]  = 0;
  ram[2913]  = 81;
  ram[2914]  = 255;
  ram[2915]  = 255;
  ram[2916]  = 255;
  ram[2917]  = 255;
  ram[2918]  = 252;
  ram[2919]  = 251;
  ram[2920]  = 238;
  ram[2921]  = 249;
  ram[2922]  = 255;
  ram[2923]  = 253;
  ram[2924]  = 253;
  ram[2925]  = 255;
  ram[2926]  = 218;
  ram[2927]  = 34;
  ram[2928]  = 0;
  ram[2929]  = 0;
  ram[2930]  = 0;
  ram[2931]  = 7;
  ram[2932]  = 1;
  ram[2933]  = 0;
  ram[2934]  = 0;
  ram[2935]  = 17;
  ram[2936]  = 182;
  ram[2937]  = 241;
  ram[2938]  = 255;
  ram[2939]  = 255;
  ram[2940]  = 255;
  ram[2941]  = 92;
  ram[2942]  = 0;
  ram[2943]  = 0;
  ram[2944]  = 3;
  ram[2945]  = 0;
  ram[2946]  = 0;
  ram[2947]  = 0;
  ram[2948]  = 0;
  ram[2949]  = 0;
  ram[2950]  = 0;
  ram[2951]  = 7;
  ram[2952]  = 0;
  ram[2953]  = 0;
  ram[2954]  = 10;
  ram[2955]  = 218;
  ram[2956]  = 255;
  ram[2957]  = 252;
  ram[2958]  = 254;
  ram[2959]  = 253;
  ram[2960]  = 255;
  ram[2961]  = 249;
  ram[2962]  = 40;
  ram[2963]  = 0;
  ram[2964]  = 0;
  ram[2965]  = 0;
  ram[2966]  = 0;
  ram[2967]  = 0;
  ram[2968]  = 0;
  ram[2969]  = 0;
  ram[2970]  = 0;
  ram[2971]  = 0;
  ram[2972]  = 13;
  ram[2973]  = 38;
  ram[2974]  = 52;
  ram[2975]  = 79;
  ram[2976]  = 106;
  ram[2977]  = 120;
  ram[2978]  = 18;
  ram[2979]  = 0;
  ram[2980]  = 0;
  ram[2981]  = 0;
  ram[2982]  = 132;
  ram[2983]  = 200;
  ram[2984]  = 222;
  ram[2985]  = 243;
  ram[2986]  = 255;
  ram[2987]  = 255;
  ram[2988]  = 255;
  ram[2989]  = 253;
  ram[2990]  = 255;
  ram[2991]  = 255;
  ram[2992]  = 255;
  ram[2993]  = 255;
  ram[2994]  = 253;
  ram[2995]  = 251;
  ram[2996]  = 252;
  ram[2997]  = 252;
  ram[2998]  = 252;
  ram[2999]  = 247;
  ram[3000]  = 244;
  ram[3001]  = 242;
  ram[3002]  = 242;
  ram[3003]  = 248;
  ram[3004]  = 243;
  ram[3005]  = 240;
  ram[3006]  = 251;
  ram[3007]  = 191;
  ram[3008]  = 81;
  ram[3009]  = 0;
  ram[3010]  = 0;
  ram[3011]  = 0;
  ram[3012]  = 0;
  ram[3013]  = 0;
  ram[3014]  = 0;
  ram[3015]  = 0;
  ram[3016]  = 125;
  ram[3017]  = 255;
  ram[3018]  = 234;
  ram[3019]  = 246;
  ram[3020]  = 214;
  ram[3021]  = 7;
  ram[3022]  = 0;
  ram[3023]  = 0;
  ram[3024]  = 168;
  ram[3025]  = 255;
  ram[3026]  = 252;
  ram[3027]  = 255;
  ram[3028]  = 255;
  ram[3029]  = 220;
  ram[3030]  = 10;
  ram[3031]  = 0;
  ram[3032]  = 0;
  ram[3033]  = 50;
  ram[3034]  = 149;
  ram[3035]  = 91;
  ram[3036]  = 62;
  ram[3037]  = 138;
  ram[3038]  = 255;
  ram[3039]  = 243;
  ram[3040]  = 231;
  ram[3041]  = 238;
  ram[3042]  = 240;
  ram[3043]  = 243;
  ram[3044]  = 242;
  ram[3045]  = 245;
  ram[3046]  = 251;
  ram[3047]  = 229;
  ram[3048]  = 150;
  ram[3049]  = 125;
  ram[3050]  = 170;
  ram[3051]  = 81;
  ram[3052]  = 0;
  ram[3053]  = 0;
  ram[3054]  = 0;
  ram[3055]  = 18;
  ram[3056]  = 182;
  ram[3057]  = 255;
  ram[3058]  = 255;
  ram[3059]  = 254;
  ram[3060]  = 255;
  ram[3061]  = 71;
  ram[3062]  = 0;
  ram[3063]  = 0;
  ram[3064]  = 0;
  ram[3065]  = 0;
  ram[3066]  = 0;
  ram[3067]  = 0;
  ram[3068]  = 0;
  ram[3069]  = 0;
  ram[3070]  = 103;
  ram[3071]  = 107;
  ram[3072]  = 0;
  ram[3073]  = 0;
  ram[3074]  = 5;
  ram[3075]  = 205;
  ram[3076]  = 252;
  ram[3077]  = 244;
  ram[3078]  = 246;
  ram[3079]  = 240;
  ram[3080]  = 243;
  ram[3081]  = 252;
  ram[3082]  = 152;
  ram[3083]  = 16;
  ram[3084]  = 0;
  ram[3085]  = 0;
  ram[3086]  = 0;
  ram[3087]  = 17;
  ram[3088]  = 56;
  ram[3089]  = 90;
  ram[3090]  = 155;
  ram[3091]  = 182;
  ram[3092]  = 220;
  ram[3093]  = 238;
  ram[3094]  = 245;
  ram[3095]  = 255;
  ram[3096]  = 255;
  ram[3097]  = 251;
  ram[3098]  = 34;
  ram[3099]  = 0;
  ram[3100]  = 0;
  ram[3101]  = 0;
  ram[3102]  = 169;
  ram[3103]  = 255;
  ram[3104]  = 253;
  ram[3105]  = 250;
  ram[3106]  = 246;
  ram[3107]  = 247;
  ram[3108]  = 238;
  ram[3109]  = 236;
  ram[3110]  = 246;
  ram[3111]  = 243;
  ram[3112]  = 239;
  ram[3113]  = 243;
  ram[3114]  = 241;
  ram[3115]  = 236;
  ram[3116]  = 240;
  ram[3117]  = 242;
  ram[3118]  = 242;
  ram[3119]  = 233;
  ram[3120]  = 244;
  ram[3121]  = 240;
  ram[3122]  = 243;
  ram[3123]  = 246;
  ram[3124]  = 243;
  ram[3125]  = 247;
  ram[3126]  = 215;
  ram[3127]  = 13;
  ram[3128]  = 0;
  ram[3129]  = 0;
  ram[3130]  = 0;
  ram[3131]  = 0;
  ram[3132]  = 0;
  ram[3133]  = 0;
  ram[3134]  = 0;
  ram[3135]  = 0;
  ram[3136]  = 121;
  ram[3137]  = 255;
  ram[3138]  = 236;
  ram[3139]  = 249;
  ram[3140]  = 203;
  ram[3141]  = 3;
  ram[3142]  = 0;
  ram[3143]  = 0;
  ram[3144]  = 177;
  ram[3145]  = 255;
  ram[3146]  = 207;
  ram[3147]  = 129;
  ram[3148]  = 76;
  ram[3149]  = 40;
  ram[3150]  = 1;
  ram[3151]  = 0;
  ram[3152]  = 0;
  ram[3153]  = 0;
  ram[3154]  = 0;
  ram[3155]  = 0;
  ram[3156]  = 0;
  ram[3157]  = 0;
  ram[3158]  = 162;
  ram[3159]  = 252;
  ram[3160]  = 237;
  ram[3161]  = 244;
  ram[3162]  = 247;
  ram[3163]  = 247;
  ram[3164]  = 246;
  ram[3165]  = 246;
  ram[3166]  = 247;
  ram[3167]  = 252;
  ram[3168]  = 255;
  ram[3169]  = 255;
  ram[3170]  = 196;
  ram[3171]  = 12;
  ram[3172]  = 0;
  ram[3173]  = 0;
  ram[3174]  = 0;
  ram[3175]  = 0;
  ram[3176]  = 0;
  ram[3177]  = 58;
  ram[3178]  = 177;
  ram[3179]  = 255;
  ram[3180]  = 253;
  ram[3181]  = 49;
  ram[3182]  = 0;
  ram[3183]  = 0;
  ram[3184]  = 17;
  ram[3185]  = 46;
  ram[3186]  = 55;
  ram[3187]  = 108;
  ram[3188]  = 171;
  ram[3189]  = 204;
  ram[3190]  = 251;
  ram[3191]  = 117;
  ram[3192]  = 0;
  ram[3193]  = 0;
  ram[3194]  = 2;
  ram[3195]  = 200;
  ram[3196]  = 255;
  ram[3197]  = 249;
  ram[3198]  = 248;
  ram[3199]  = 246;
  ram[3200]  = 246;
  ram[3201]  = 249;
  ram[3202]  = 255;
  ram[3203]  = 216;
  ram[3204]  = 154;
  ram[3205]  = 156;
  ram[3206]  = 184;
  ram[3207]  = 227;
  ram[3208]  = 255;
  ram[3209]  = 255;
  ram[3210]  = 255;
  ram[3211]  = 255;
  ram[3212]  = 255;
  ram[3213]  = 253;
  ram[3214]  = 248;
  ram[3215]  = 251;
  ram[3216]  = 253;
  ram[3217]  = 240;
  ram[3218]  = 41;
  ram[3219]  = 0;
  ram[3220]  = 0;
  ram[3221]  = 0;
  ram[3222]  = 130;
  ram[3223]  = 255;
  ram[3224]  = 250;
  ram[3225]  = 250;
  ram[3226]  = 249;
  ram[3227]  = 251;
  ram[3228]  = 241;
  ram[3229]  = 240;
  ram[3230]  = 249;
  ram[3231]  = 247;
  ram[3232]  = 245;
  ram[3233]  = 249;
  ram[3234]  = 248;
  ram[3235]  = 247;
  ram[3236]  = 249;
  ram[3237]  = 249;
  ram[3238]  = 248;
  ram[3239]  = 241;
  ram[3240]  = 251;
  ram[3241]  = 253;
  ram[3242]  = 253;
  ram[3243]  = 252;
  ram[3244]  = 254;
  ram[3245]  = 255;
  ram[3246]  = 202;
  ram[3247]  = 0;
  ram[3248]  = 0;
  ram[3249]  = 0;
  ram[3250]  = 0;
  ram[3251]  = 37;
  ram[3252]  = 124;
  ram[3253]  = 11;
  ram[3254]  = 0;
  ram[3255]  = 0;
  ram[3256]  = 119;
  ram[3257]  = 255;
  ram[3258]  = 244;
  ram[3259]  = 255;
  ram[3260]  = 200;
  ram[3261]  = 0;
  ram[3262]  = 0;
  ram[3263]  = 0;
  ram[3264]  = 201;
  ram[3265]  = 193;
  ram[3266]  = 8;
  ram[3267]  = 0;
  ram[3268]  = 0;
  ram[3269]  = 0;
  ram[3270]  = 0;
  ram[3271]  = 0;
  ram[3272]  = 0;
  ram[3273]  = 0;
  ram[3274]  = 0;
  ram[3275]  = 0;
  ram[3276]  = 0;
  ram[3277]  = 0;
  ram[3278]  = 137;
  ram[3279]  = 255;
  ram[3280]  = 242;
  ram[3281]  = 250;
  ram[3282]  = 255;
  ram[3283]  = 254;
  ram[3284]  = 254;
  ram[3285]  = 254;
  ram[3286]  = 253;
  ram[3287]  = 252;
  ram[3288]  = 255;
  ram[3289]  = 218;
  ram[3290]  = 27;
  ram[3291]  = 0;
  ram[3292]  = 0;
  ram[3293]  = 0;
  ram[3294]  = 0;
  ram[3295]  = 0;
  ram[3296]  = 0;
  ram[3297]  = 0;
  ram[3298]  = 0;
  ram[3299]  = 126;
  ram[3300]  = 255;
  ram[3301]  = 62;
  ram[3302]  = 0;
  ram[3303]  = 0;
  ram[3304]  = 76;
  ram[3305]  = 255;
  ram[3306]  = 255;
  ram[3307]  = 255;
  ram[3308]  = 255;
  ram[3309]  = 255;
  ram[3310]  = 255;
  ram[3311]  = 117;
  ram[3312]  = 0;
  ram[3313]  = 0;
  ram[3314]  = 0;
  ram[3315]  = 186;
  ram[3316]  = 255;
  ram[3317]  = 253;
  ram[3318]  = 252;
  ram[3319]  = 251;
  ram[3320]  = 254;
  ram[3321]  = 252;
  ram[3322]  = 253;
  ram[3323]  = 255;
  ram[3324]  = 255;
  ram[3325]  = 255;
  ram[3326]  = 255;
  ram[3327]  = 255;
  ram[3328]  = 255;
  ram[3329]  = 254;
  ram[3330]  = 253;
  ram[3331]  = 253;
  ram[3332]  = 254;
  ram[3333]  = 253;
  ram[3334]  = 252;
  ram[3335]  = 253;
  ram[3336]  = 255;
  ram[3337]  = 249;
  ram[3338]  = 50;
  ram[3339]  = 0;
  ram[3340]  = 0;
  ram[3341]  = 0;
  ram[3342]  = 115;
  ram[3343]  = 255;
  ram[3344]  = 254;
  ram[3345]  = 253;
  ram[3346]  = 254;
  ram[3347]  = 254;
  ram[3348]  = 245;
  ram[3349]  = 244;
  ram[3350]  = 253;
  ram[3351]  = 251;
  ram[3352]  = 250;
  ram[3353]  = 252;
  ram[3354]  = 253;
  ram[3355]  = 252;
  ram[3356]  = 253;
  ram[3357]  = 252;
  ram[3358]  = 252;
  ram[3359]  = 247;
  ram[3360]  = 251;
  ram[3361]  = 252;
  ram[3362]  = 253;
  ram[3363]  = 253;
  ram[3364]  = 253;
  ram[3365]  = 255;
  ram[3366]  = 251;
  ram[3367]  = 89;
  ram[3368]  = 0;
  ram[3369]  = 3;
  ram[3370]  = 108;
  ram[3371]  = 241;
  ram[3372]  = 225;
  ram[3373]  = 6;
  ram[3374]  = 0;
  ram[3375]  = 0;
  ram[3376]  = 114;
  ram[3377]  = 255;
  ram[3378]  = 245;
  ram[3379]  = 254;
  ram[3380]  = 202;
  ram[3381]  = 0;
  ram[3382]  = 0;
  ram[3383]  = 0;
  ram[3384]  = 190;
  ram[3385]  = 192;
  ram[3386]  = 0;
  ram[3387]  = 0;
  ram[3388]  = 0;
  ram[3389]  = 0;
  ram[3390]  = 0;
  ram[3391]  = 0;
  ram[3392]  = 0;
  ram[3393]  = 8;
  ram[3394]  = 49;
  ram[3395]  = 90;
  ram[3396]  = 110;
  ram[3397]  = 199;
  ram[3398]  = 251;
  ram[3399]  = 252;
  ram[3400]  = 242;
  ram[3401]  = 249;
  ram[3402]  = 254;
  ram[3403]  = 253;
  ram[3404]  = 253;
  ram[3405]  = 252;
  ram[3406]  = 252;
  ram[3407]  = 255;
  ram[3408]  = 255;
  ram[3409]  = 69;
  ram[3410]  = 0;
  ram[3411]  = 0;
  ram[3412]  = 0;
  ram[3413]  = 0;
  ram[3414]  = 0;
  ram[3415]  = 8;
  ram[3416]  = 4;
  ram[3417]  = 0;
  ram[3418]  = 0;
  ram[3419]  = 0;
  ram[3420]  = 175;
  ram[3421]  = 99;
  ram[3422]  = 0;
  ram[3423]  = 0;
  ram[3424]  = 65;
  ram[3425]  = 255;
  ram[3426]  = 243;
  ram[3427]  = 203;
  ram[3428]  = 174;
  ram[3429]  = 154;
  ram[3430]  = 150;
  ram[3431]  = 78;
  ram[3432]  = 0;
  ram[3433]  = 0;
  ram[3434]  = 0;
  ram[3435]  = 176;
  ram[3436]  = 255;
  ram[3437]  = 252;
  ram[3438]  = 252;
  ram[3439]  = 252;
  ram[3440]  = 253;
  ram[3441]  = 250;
  ram[3442]  = 252;
  ram[3443]  = 253;
  ram[3444]  = 253;
  ram[3445]  = 249;
  ram[3446]  = 242;
  ram[3447]  = 252;
  ram[3448]  = 253;
  ram[3449]  = 253;
  ram[3450]  = 253;
  ram[3451]  = 252;
  ram[3452]  = 252;
  ram[3453]  = 253;
  ram[3454]  = 252;
  ram[3455]  = 253;
  ram[3456]  = 255;
  ram[3457]  = 247;
  ram[3458]  = 45;
  ram[3459]  = 0;
  ram[3460]  = 0;
  ram[3461]  = 0;
  ram[3462]  = 108;
  ram[3463]  = 255;
  ram[3464]  = 253;
  ram[3465]  = 252;
  ram[3466]  = 253;
  ram[3467]  = 253;
  ram[3468]  = 244;
  ram[3469]  = 244;
  ram[3470]  = 252;
  ram[3471]  = 250;
  ram[3472]  = 250;
  ram[3473]  = 250;
  ram[3474]  = 252;
  ram[3475]  = 251;
  ram[3476]  = 250;
  ram[3477]  = 251;
  ram[3478]  = 251;
  ram[3479]  = 242;
  ram[3480]  = 251;
  ram[3481]  = 251;
  ram[3482]  = 251;
  ram[3483]  = 252;
  ram[3484]  = 254;
  ram[3485]  = 253;
  ram[3486]  = 255;
  ram[3487]  = 255;
  ram[3488]  = 200;
  ram[3489]  = 198;
  ram[3490]  = 255;
  ram[3491]  = 255;
  ram[3492]  = 201;
  ram[3493]  = 1;
  ram[3494]  = 0;
  ram[3495]  = 0;
  ram[3496]  = 112;
  ram[3497]  = 255;
  ram[3498]  = 245;
  ram[3499]  = 253;
  ram[3500]  = 207;
  ram[3501]  = 3;
  ram[3502]  = 0;
  ram[3503]  = 0;
  ram[3504]  = 173;
  ram[3505]  = 255;
  ram[3506]  = 154;
  ram[3507]  = 58;
  ram[3508]  = 60;
  ram[3509]  = 95;
  ram[3510]  = 19;
  ram[3511]  = 0;
  ram[3512]  = 0;
  ram[3513]  = 73;
  ram[3514]  = 254;
  ram[3515]  = 255;
  ram[3516]  = 255;
  ram[3517]  = 255;
  ram[3518]  = 254;
  ram[3519]  = 251;
  ram[3520]  = 244;
  ram[3521]  = 251;
  ram[3522]  = 253;
  ram[3523]  = 253;
  ram[3524]  = 252;
  ram[3525]  = 252;
  ram[3526]  = 253;
  ram[3527]  = 255;
  ram[3528]  = 116;
  ram[3529]  = 0;
  ram[3530]  = 0;
  ram[3531]  = 0;
  ram[3532]  = 10;
  ram[3533]  = 2;
  ram[3534]  = 0;
  ram[3535]  = 26;
  ram[3536]  = 161;
  ram[3537]  = 22;
  ram[3538]  = 0;
  ram[3539]  = 0;
  ram[3540]  = 134;
  ram[3541]  = 99;
  ram[3542]  = 0;
  ram[3543]  = 0;
  ram[3544]  = 25;
  ram[3545]  = 64;
  ram[3546]  = 26;
  ram[3547]  = 0;
  ram[3548]  = 0;
  ram[3549]  = 0;
  ram[3550]  = 0;
  ram[3551]  = 0;
  ram[3552]  = 0;
  ram[3553]  = 0;
  ram[3554]  = 0;
  ram[3555]  = 189;
  ram[3556]  = 255;
  ram[3557]  = 252;
  ram[3558]  = 252;
  ram[3559]  = 250;
  ram[3560]  = 252;
  ram[3561]  = 251;
  ram[3562]  = 253;
  ram[3563]  = 252;
  ram[3564]  = 253;
  ram[3565]  = 248;
  ram[3566]  = 244;
  ram[3567]  = 252;
  ram[3568]  = 253;
  ram[3569]  = 251;
  ram[3570]  = 251;
  ram[3571]  = 252;
  ram[3572]  = 252;
  ram[3573]  = 253;
  ram[3574]  = 253;
  ram[3575]  = 253;
  ram[3576]  = 254;
  ram[3577]  = 249;
  ram[3578]  = 49;
  ram[3579]  = 0;
  ram[3580]  = 0;
  ram[3581]  = 0;
  ram[3582]  = 112;
  ram[3583]  = 255;
  ram[3584]  = 253;
  ram[3585]  = 251;
  ram[3586]  = 252;
  ram[3587]  = 253;
  ram[3588]  = 245;
  ram[3589]  = 244;
  ram[3590]  = 253;
  ram[3591]  = 251;
  ram[3592]  = 251;
  ram[3593]  = 251;
  ram[3594]  = 251;
  ram[3595]  = 251;
  ram[3596]  = 249;
  ram[3597]  = 250;
  ram[3598]  = 251;
  ram[3599]  = 245;
  ram[3600]  = 251;
  ram[3601]  = 251;
  ram[3602]  = 252;
  ram[3603]  = 252;
  ram[3604]  = 253;
  ram[3605]  = 253;
  ram[3606]  = 252;
  ram[3607]  = 255;
  ram[3608]  = 255;
  ram[3609]  = 253;
  ram[3610]  = 253;
  ram[3611]  = 255;
  ram[3612]  = 200;
  ram[3613]  = 1;
  ram[3614]  = 0;
  ram[3615]  = 0;
  ram[3616]  = 116;
  ram[3617]  = 255;
  ram[3618]  = 243;
  ram[3619]  = 254;
  ram[3620]  = 208;
  ram[3621]  = 7;
  ram[3622]  = 0;
  ram[3623]  = 0;
  ram[3624]  = 151;
  ram[3625]  = 255;
  ram[3626]  = 255;
  ram[3627]  = 255;
  ram[3628]  = 255;
  ram[3629]  = 242;
  ram[3630]  = 20;
  ram[3631]  = 0;
  ram[3632]  = 0;
  ram[3633]  = 86;
  ram[3634]  = 255;
  ram[3635]  = 255;
  ram[3636]  = 255;
  ram[3637]  = 255;
  ram[3638]  = 255;
  ram[3639]  = 255;
  ram[3640]  = 246;
  ram[3641]  = 251;
  ram[3642]  = 253;
  ram[3643]  = 252;
  ram[3644]  = 252;
  ram[3645]  = 252;
  ram[3646]  = 255;
  ram[3647]  = 160;
  ram[3648]  = 0;
  ram[3649]  = 0;
  ram[3650]  = 0;
  ram[3651]  = 32;
  ram[3652]  = 111;
  ram[3653]  = 0;
  ram[3654]  = 0;
  ram[3655]  = 20;
  ram[3656]  = 248;
  ram[3657]  = 213;
  ram[3658]  = 70;
  ram[3659]  = 85;
  ram[3660]  = 242;
  ram[3661]  = 73;
  ram[3662]  = 0;
  ram[3663]  = 0;
  ram[3664]  = 0;
  ram[3665]  = 0;
  ram[3666]  = 0;
  ram[3667]  = 0;
  ram[3668]  = 0;
  ram[3669]  = 0;
  ram[3670]  = 5;
  ram[3671]  = 15;
  ram[3672]  = 0;
  ram[3673]  = 0;
  ram[3674]  = 0;
  ram[3675]  = 185;
  ram[3676]  = 255;
  ram[3677]  = 252;
  ram[3678]  = 251;
  ram[3679]  = 250;
  ram[3680]  = 252;
  ram[3681]  = 252;
  ram[3682]  = 252;
  ram[3683]  = 252;
  ram[3684]  = 251;
  ram[3685]  = 247;
  ram[3686]  = 246;
  ram[3687]  = 253;
  ram[3688]  = 252;
  ram[3689]  = 250;
  ram[3690]  = 250;
  ram[3691]  = 252;
  ram[3692]  = 252;
  ram[3693]  = 253;
  ram[3694]  = 253;
  ram[3695]  = 252;
  ram[3696]  = 255;
  ram[3697]  = 235;
  ram[3698]  = 28;
  ram[3699]  = 0;
  ram[3700]  = 0;
  ram[3701]  = 0;
  ram[3702]  = 115;
  ram[3703]  = 255;
  ram[3704]  = 253;
  ram[3705]  = 251;
  ram[3706]  = 250;
  ram[3707]  = 253;
  ram[3708]  = 247;
  ram[3709]  = 245;
  ram[3710]  = 252;
  ram[3711]  = 251;
  ram[3712]  = 252;
  ram[3713]  = 251;
  ram[3714]  = 249;
  ram[3715]  = 251;
  ram[3716]  = 251;
  ram[3717]  = 250;
  ram[3718]  = 252;
  ram[3719]  = 245;
  ram[3720]  = 252;
  ram[3721]  = 252;
  ram[3722]  = 251;
  ram[3723]  = 252;
  ram[3724]  = 251;
  ram[3725]  = 252;
  ram[3726]  = 253;
  ram[3727]  = 252;
  ram[3728]  = 249;
  ram[3729]  = 253;
  ram[3730]  = 255;
  ram[3731]  = 255;
  ram[3732]  = 195;
  ram[3733]  = 0;
  ram[3734]  = 0;
  ram[3735]  = 0;
  ram[3736]  = 133;
  ram[3737]  = 255;
  ram[3738]  = 245;
  ram[3739]  = 255;
  ram[3740]  = 183;
  ram[3741]  = 0;
  ram[3742]  = 0;
  ram[3743]  = 0;
  ram[3744]  = 166;
  ram[3745]  = 255;
  ram[3746]  = 252;
  ram[3747]  = 255;
  ram[3748]  = 255;
  ram[3749]  = 247;
  ram[3750]  = 31;
  ram[3751]  = 0;
  ram[3752]  = 0;
  ram[3753]  = 98;
  ram[3754]  = 255;
  ram[3755]  = 255;
  ram[3756]  = 255;
  ram[3757]  = 255;
  ram[3758]  = 254;
  ram[3759]  = 244;
  ram[3760]  = 255;
  ram[3761]  = 255;
  ram[3762]  = 252;
  ram[3763]  = 252;
  ram[3764]  = 253;
  ram[3765]  = 255;
  ram[3766]  = 202;
  ram[3767]  = 13;
  ram[3768]  = 0;
  ram[3769]  = 0;
  ram[3770]  = 0;
  ram[3771]  = 171;
  ram[3772]  = 149;
  ram[3773]  = 0;
  ram[3774]  = 0;
  ram[3775]  = 18;
  ram[3776]  = 227;
  ram[3777]  = 255;
  ram[3778]  = 255;
  ram[3779]  = 255;
  ram[3780]  = 255;
  ram[3781]  = 55;
  ram[3782]  = 0;
  ram[3783]  = 0;
  ram[3784]  = 0;
  ram[3785]  = 0;
  ram[3786]  = 14;
  ram[3787]  = 48;
  ram[3788]  = 80;
  ram[3789]  = 100;
  ram[3790]  = 194;
  ram[3791]  = 98;
  ram[3792]  = 0;
  ram[3793]  = 0;
  ram[3794]  = 0;
  ram[3795]  = 173;
  ram[3796]  = 255;
  ram[3797]  = 253;
  ram[3798]  = 251;
  ram[3799]  = 250;
  ram[3800]  = 251;
  ram[3801]  = 252;
  ram[3802]  = 252;
  ram[3803]  = 253;
  ram[3804]  = 254;
  ram[3805]  = 247;
  ram[3806]  = 242;
  ram[3807]  = 253;
  ram[3808]  = 252;
  ram[3809]  = 253;
  ram[3810]  = 253;
  ram[3811]  = 252;
  ram[3812]  = 251;
  ram[3813]  = 252;
  ram[3814]  = 252;
  ram[3815]  = 253;
  ram[3816]  = 255;
  ram[3817]  = 218;
  ram[3818]  = 6;
  ram[3819]  = 0;
  ram[3820]  = 0;
  ram[3821]  = 0;
  ram[3822]  = 146;
  ram[3823]  = 255;
  ram[3824]  = 252;
  ram[3825]  = 251;
  ram[3826]  = 252;
  ram[3827]  = 254;
  ram[3828]  = 244;
  ram[3829]  = 241;
  ram[3830]  = 251;
  ram[3831]  = 252;
  ram[3832]  = 252;
  ram[3833]  = 250;
  ram[3834]  = 250;
  ram[3835]  = 251;
  ram[3836]  = 250;
  ram[3837]  = 251;
  ram[3838]  = 253;
  ram[3839]  = 241;
  ram[3840]  = 252;
  ram[3841]  = 251;
  ram[3842]  = 252;
  ram[3843]  = 251;
  ram[3844]  = 251;
  ram[3845]  = 252;
  ram[3846]  = 252;
  ram[3847]  = 253;
  ram[3848]  = 246;
  ram[3849]  = 198;
  ram[3850]  = 253;
  ram[3851]  = 255;
  ram[3852]  = 169;
  ram[3853]  = 0;
  ram[3854]  = 0;
  ram[3855]  = 0;
  ram[3856]  = 156;
  ram[3857]  = 255;
  ram[3858]  = 246;
  ram[3859]  = 255;
  ram[3860]  = 179;
  ram[3861]  = 0;
  ram[3862]  = 0;
  ram[3863]  = 0;
  ram[3864]  = 167;
  ram[3865]  = 255;
  ram[3866]  = 255;
  ram[3867]  = 255;
  ram[3868]  = 246;
  ram[3869]  = 191;
  ram[3870]  = 11;
  ram[3871]  = 0;
  ram[3872]  = 0;
  ram[3873]  = 36;
  ram[3874]  = 90;
  ram[3875]  = 76;
  ram[3876]  = 67;
  ram[3877]  = 52;
  ram[3878]  = 51;
  ram[3879]  = 35;
  ram[3880]  = 110;
  ram[3881]  = 232;
  ram[3882]  = 255;
  ram[3883]  = 253;
  ram[3884]  = 254;
  ram[3885]  = 250;
  ram[3886]  = 59;
  ram[3887]  = 0;
  ram[3888]  = 0;
  ram[3889]  = 0;
  ram[3890]  = 90;
  ram[3891]  = 255;
  ram[3892]  = 140;
  ram[3893]  = 0;
  ram[3894]  = 0;
  ram[3895]  = 19;
  ram[3896]  = 229;
  ram[3897]  = 255;
  ram[3898]  = 253;
  ram[3899]  = 255;
  ram[3900]  = 251;
  ram[3901]  = 48;
  ram[3902]  = 0;
  ram[3903]  = 0;
  ram[3904]  = 46;
  ram[3905]  = 200;
  ram[3906]  = 225;
  ram[3907]  = 255;
  ram[3908]  = 255;
  ram[3909]  = 255;
  ram[3910]  = 255;
  ram[3911]  = 92;
  ram[3912]  = 0;
  ram[3913]  = 0;
  ram[3914]  = 8;
  ram[3915]  = 177;
  ram[3916]  = 255;
  ram[3917]  = 252;
  ram[3918]  = 251;
  ram[3919]  = 252;
  ram[3920]  = 252;
  ram[3921]  = 252;
  ram[3922]  = 253;
  ram[3923]  = 252;
  ram[3924]  = 254;
  ram[3925]  = 249;
  ram[3926]  = 242;
  ram[3927]  = 252;
  ram[3928]  = 252;
  ram[3929]  = 252;
  ram[3930]  = 253;
  ram[3931]  = 252;
  ram[3932]  = 255;
  ram[3933]  = 255;
  ram[3934]  = 255;
  ram[3935]  = 254;
  ram[3936]  = 255;
  ram[3937]  = 192;
  ram[3938]  = 0;
  ram[3939]  = 0;
  ram[3940]  = 0;
  ram[3941]  = 0;
  ram[3942]  = 177;
  ram[3943]  = 255;
  ram[3944]  = 252;
  ram[3945]  = 252;
  ram[3946]  = 252;
  ram[3947]  = 253;
  ram[3948]  = 245;
  ram[3949]  = 243;
  ram[3950]  = 251;
  ram[3951]  = 251;
  ram[3952]  = 251;
  ram[3953]  = 250;
  ram[3954]  = 251;
  ram[3955]  = 250;
  ram[3956]  = 250;
  ram[3957]  = 252;
  ram[3958]  = 253;
  ram[3959]  = 244;
  ram[3960]  = 251;
  ram[3961]  = 250;
  ram[3962]  = 252;
  ram[3963]  = 251;
  ram[3964]  = 251;
  ram[3965]  = 253;
  ram[3966]  = 252;
  ram[3967]  = 255;
  ram[3968]  = 230;
  ram[3969]  = 73;
  ram[3970]  = 65;
  ram[3971]  = 159;
  ram[3972]  = 97;
  ram[3973]  = 0;
  ram[3974]  = 0;
  ram[3975]  = 0;
  ram[3976]  = 180;
  ram[3977]  = 255;
  ram[3978]  = 246;
  ram[3979]  = 255;
  ram[3980]  = 178;
  ram[3981]  = 0;
  ram[3982]  = 0;
  ram[3983]  = 0;
  ram[3984]  = 164;
  ram[3985]  = 168;
  ram[3986]  = 97;
  ram[3987]  = 68;
  ram[3988]  = 35;
  ram[3989]  = 2;
  ram[3990]  = 0;
  ram[3991]  = 0;
  ram[3992]  = 0;
  ram[3993]  = 0;
  ram[3994]  = 0;
  ram[3995]  = 0;
  ram[3996]  = 0;
  ram[3997]  = 0;
  ram[3998]  = 0;
  ram[3999]  = 0;
  ram[4000]  = 0;
  ram[4001]  = 60;
  ram[4002]  = 246;
  ram[4003]  = 255;
  ram[4004]  = 255;
  ram[4005]  = 248;
  ram[4006]  = 44;
  ram[4007]  = 0;
  ram[4008]  = 0;
  ram[4009]  = 68;
  ram[4010]  = 238;
  ram[4011]  = 255;
  ram[4012]  = 131;
  ram[4013]  = 0;
  ram[4014]  = 0;
  ram[4015]  = 18;
  ram[4016]  = 228;
  ram[4017]  = 255;
  ram[4018]  = 251;
  ram[4019]  = 255;
  ram[4020]  = 239;
  ram[4021]  = 27;
  ram[4022]  = 0;
  ram[4023]  = 0;
  ram[4024]  = 48;
  ram[4025]  = 255;
  ram[4026]  = 255;
  ram[4027]  = 255;
  ram[4028]  = 255;
  ram[4029]  = 255;
  ram[4030]  = 247;
  ram[4031]  = 59;
  ram[4032]  = 0;
  ram[4033]  = 1;
  ram[4034]  = 10;
  ram[4035]  = 185;
  ram[4036]  = 255;
  ram[4037]  = 252;
  ram[4038]  = 251;
  ram[4039]  = 251;
  ram[4040]  = 253;
  ram[4041]  = 252;
  ram[4042]  = 253;
  ram[4043]  = 253;
  ram[4044]  = 254;
  ram[4045]  = 248;
  ram[4046]  = 242;
  ram[4047]  = 252;
  ram[4048]  = 253;
  ram[4049]  = 252;
  ram[4050]  = 252;
  ram[4051]  = 251;
  ram[4052]  = 234;
  ram[4053]  = 210;
  ram[4054]  = 241;
  ram[4055]  = 255;
  ram[4056]  = 255;
  ram[4057]  = 126;
  ram[4058]  = 0;
  ram[4059]  = 0;
  ram[4060]  = 0;
  ram[4061]  = 0;
  ram[4062]  = 200;
  ram[4063]  = 255;
  ram[4064]  = 252;
  ram[4065]  = 251;
  ram[4066]  = 251;
  ram[4067]  = 252;
  ram[4068]  = 245;
  ram[4069]  = 245;
  ram[4070]  = 253;
  ram[4071]  = 251;
  ram[4072]  = 251;
  ram[4073]  = 250;
  ram[4074]  = 250;
  ram[4075]  = 251;
  ram[4076]  = 252;
  ram[4077]  = 252;
  ram[4078]  = 253;
  ram[4079]  = 244;
  ram[4080]  = 251;
  ram[4081]  = 251;
  ram[4082]  = 252;
  ram[4083]  = 251;
  ram[4084]  = 250;
  ram[4085]  = 251;
  ram[4086]  = 251;
  ram[4087]  = 253;
  ram[4088]  = 249;
  ram[4089]  = 116;
  ram[4090]  = 0;
  ram[4091]  = 0;
  ram[4092]  = 0;
  ram[4093]  = 0;
  ram[4094]  = 0;
  ram[4095]  = 12;
  ram[4096]  = 225;
  ram[4097]  = 255;
  ram[4098]  = 246;
  ram[4099]  = 255;
  ram[4100]  = 160;
  ram[4101]  = 0;
  ram[4102]  = 0;
  ram[4103]  = 1;
  ram[4104]  = 44;
  ram[4105]  = 0;
  ram[4106]  = 0;
  ram[4107]  = 0;
  ram[4108]  = 0;
  ram[4109]  = 0;
  ram[4110]  = 0;
  ram[4111]  = 0;
  ram[4112]  = 0;
  ram[4113]  = 0;
  ram[4114]  = 0;
  ram[4115]  = 0;
  ram[4116]  = 0;
  ram[4117]  = 0;
  ram[4118]  = 0;
  ram[4119]  = 0;
  ram[4120]  = 0;
  ram[4121]  = 33;
  ram[4122]  = 242;
  ram[4123]  = 255;
  ram[4124]  = 253;
  ram[4125]  = 254;
  ram[4126]  = 205;
  ram[4127]  = 67;
  ram[4128]  = 85;
  ram[4129]  = 245;
  ram[4130]  = 255;
  ram[4131]  = 255;
  ram[4132]  = 106;
  ram[4133]  = 0;
  ram[4134]  = 0;
  ram[4135]  = 9;
  ram[4136]  = 217;
  ram[4137]  = 255;
  ram[4138]  = 251;
  ram[4139]  = 254;
  ram[4140]  = 243;
  ram[4141]  = 42;
  ram[4142]  = 0;
  ram[4143]  = 0;
  ram[4144]  = 25;
  ram[4145]  = 180;
  ram[4146]  = 151;
  ram[4147]  = 97;
  ram[4148]  = 87;
  ram[4149]  = 65;
  ram[4150]  = 39;
  ram[4151]  = 6;
  ram[4152]  = 0;
  ram[4153]  = 3;
  ram[4154]  = 25;
  ram[4155]  = 187;
  ram[4156]  = 255;
  ram[4157]  = 252;
  ram[4158]  = 251;
  ram[4159]  = 252;
  ram[4160]  = 252;
  ram[4161]  = 253;
  ram[4162]  = 252;
  ram[4163]  = 253;
  ram[4164]  = 253;
  ram[4165]  = 247;
  ram[4166]  = 241;
  ram[4167]  = 251;
  ram[4168]  = 253;
  ram[4169]  = 253;
  ram[4170]  = 254;
  ram[4171]  = 251;
  ram[4172]  = 150;
  ram[4173]  = 80;
  ram[4174]  = 67;
  ram[4175]  = 134;
  ram[4176]  = 156;
  ram[4177]  = 18;
  ram[4178]  = 0;
  ram[4179]  = 0;
  ram[4180]  = 0;
  ram[4181]  = 51;
  ram[4182]  = 245;
  ram[4183]  = 255;
  ram[4184]  = 252;
  ram[4185]  = 251;
  ram[4186]  = 250;
  ram[4187]  = 251;
  ram[4188]  = 243;
  ram[4189]  = 245;
  ram[4190]  = 253;
  ram[4191]  = 251;
  ram[4192]  = 251;
  ram[4193]  = 251;
  ram[4194]  = 250;
  ram[4195]  = 250;
  ram[4196]  = 253;
  ram[4197]  = 253;
  ram[4198]  = 253;
  ram[4199]  = 243;
  ram[4200]  = 252;
  ram[4201]  = 251;
  ram[4202]  = 251;
  ram[4203]  = 252;
  ram[4204]  = 251;
  ram[4205]  = 250;
  ram[4206]  = 250;
  ram[4207]  = 251;
  ram[4208]  = 255;
  ram[4209]  = 218;
  ram[4210]  = 40;
  ram[4211]  = 0;
  ram[4212]  = 0;
  ram[4213]  = 0;
  ram[4214]  = 0;
  ram[4215]  = 46;
  ram[4216]  = 250;
  ram[4217]  = 255;
  ram[4218]  = 245;
  ram[4219]  = 255;
  ram[4220]  = 154;
  ram[4221]  = 0;
  ram[4222]  = 0;
  ram[4223]  = 0;
  ram[4224]  = 0;
  ram[4225]  = 0;
  ram[4226]  = 0;
  ram[4227]  = 0;
  ram[4228]  = 0;
  ram[4229]  = 0;
  ram[4230]  = 0;
  ram[4231]  = 0;
  ram[4232]  = 0;
  ram[4233]  = 26;
  ram[4234]  = 35;
  ram[4235]  = 38;
  ram[4236]  = 37;
  ram[4237]  = 19;
  ram[4238]  = 3;
  ram[4239]  = 21;
  ram[4240]  = 56;
  ram[4241]  = 183;
  ram[4242]  = 255;
  ram[4243]  = 252;
  ram[4244]  = 252;
  ram[4245]  = 251;
  ram[4246]  = 255;
  ram[4247]  = 253;
  ram[4248]  = 255;
  ram[4249]  = 255;
  ram[4250]  = 254;
  ram[4251]  = 255;
  ram[4252]  = 90;
  ram[4253]  = 0;
  ram[4254]  = 0;
  ram[4255]  = 15;
  ram[4256]  = 224;
  ram[4257]  = 255;
  ram[4258]  = 251;
  ram[4259]  = 253;
  ram[4260]  = 255;
  ram[4261]  = 93;
  ram[4262]  = 0;
  ram[4263]  = 0;
  ram[4264]  = 0;
  ram[4265]  = 0;
  ram[4266]  = 0;
  ram[4267]  = 0;
  ram[4268]  = 0;
  ram[4269]  = 0;
  ram[4270]  = 0;
  ram[4271]  = 0;
  ram[4272]  = 0;
  ram[4273]  = 0;
  ram[4274]  = 11;
  ram[4275]  = 209;
  ram[4276]  = 255;
  ram[4277]  = 252;
  ram[4278]  = 252;
  ram[4279]  = 253;
  ram[4280]  = 252;
  ram[4281]  = 252;
  ram[4282]  = 252;
  ram[4283]  = 252;
  ram[4284]  = 253;
  ram[4285]  = 247;
  ram[4286]  = 241;
  ram[4287]  = 252;
  ram[4288]  = 253;
  ram[4289]  = 253;
  ram[4290]  = 253;
  ram[4291]  = 255;
  ram[4292]  = 189;
  ram[4293]  = 11;
  ram[4294]  = 0;
  ram[4295]  = 0;
  ram[4296]  = 0;
  ram[4297]  = 0;
  ram[4298]  = 0;
  ram[4299]  = 0;
  ram[4300]  = 0;
  ram[4301]  = 121;
  ram[4302]  = 255;
  ram[4303]  = 252;
  ram[4304]  = 253;
  ram[4305]  = 251;
  ram[4306]  = 249;
  ram[4307]  = 251;
  ram[4308]  = 242;
  ram[4309]  = 243;
  ram[4310]  = 251;
  ram[4311]  = 250;
  ram[4312]  = 251;
  ram[4313]  = 251;
  ram[4314]  = 250;
  ram[4315]  = 251;
  ram[4316]  = 252;
  ram[4317]  = 253;
  ram[4318]  = 253;
  ram[4319]  = 243;
  ram[4320]  = 254;
  ram[4321]  = 253;
  ram[4322]  = 254;
  ram[4323]  = 252;
  ram[4324]  = 251;
  ram[4325]  = 250;
  ram[4326]  = 250;
  ram[4327]  = 251;
  ram[4328]  = 251;
  ram[4329]  = 255;
  ram[4330]  = 134;
  ram[4331]  = 0;
  ram[4332]  = 0;
  ram[4333]  = 0;
  ram[4334]  = 0;
  ram[4335]  = 120;
  ram[4336]  = 255;
  ram[4337]  = 254;
  ram[4338]  = 245;
  ram[4339]  = 255;
  ram[4340]  = 162;
  ram[4341]  = 0;
  ram[4342]  = 0;
  ram[4343]  = 0;
  ram[4344]  = 103;
  ram[4345]  = 130;
  ram[4346]  = 66;
  ram[4347]  = 64;
  ram[4348]  = 101;
  ram[4349]  = 110;
  ram[4350]  = 142;
  ram[4351]  = 162;
  ram[4352]  = 197;
  ram[4353]  = 235;
  ram[4354]  = 244;
  ram[4355]  = 246;
  ram[4356]  = 246;
  ram[4357]  = 231;
  ram[4358]  = 212;
  ram[4359]  = 228;
  ram[4360]  = 249;
  ram[4361]  = 255;
  ram[4362]  = 254;
  ram[4363]  = 253;
  ram[4364]  = 253;
  ram[4365]  = 252;
  ram[4366]  = 251;
  ram[4367]  = 255;
  ram[4368]  = 255;
  ram[4369]  = 253;
  ram[4370]  = 254;
  ram[4371]  = 255;
  ram[4372]  = 95;
  ram[4373]  = 0;
  ram[4374]  = 0;
  ram[4375]  = 5;
  ram[4376]  = 215;
  ram[4377]  = 255;
  ram[4378]  = 251;
  ram[4379]  = 252;
  ram[4380]  = 255;
  ram[4381]  = 168;
  ram[4382]  = 0;
  ram[4383]  = 0;
  ram[4384]  = 0;
  ram[4385]  = 0;
  ram[4386]  = 0;
  ram[4387]  = 0;
  ram[4388]  = 0;
  ram[4389]  = 0;
  ram[4390]  = 0;
  ram[4391]  = 0;
  ram[4392]  = 0;
  ram[4393]  = 0;
  ram[4394]  = 11;
  ram[4395]  = 216;
  ram[4396]  = 255;
  ram[4397]  = 252;
  ram[4398]  = 251;
  ram[4399]  = 252;
  ram[4400]  = 252;
  ram[4401]  = 253;
  ram[4402]  = 253;
  ram[4403]  = 252;
  ram[4404]  = 254;
  ram[4405]  = 248;
  ram[4406]  = 241;
  ram[4407]  = 253;
  ram[4408]  = 253;
  ram[4409]  = 253;
  ram[4410]  = 252;
  ram[4411]  = 254;
  ram[4412]  = 247;
  ram[4413]  = 57;
  ram[4414]  = 0;
  ram[4415]  = 0;
  ram[4416]  = 0;
  ram[4417]  = 0;
  ram[4418]  = 0;
  ram[4419]  = 0;
  ram[4420]  = 12;
  ram[4421]  = 210;
  ram[4422]  = 255;
  ram[4423]  = 251;
  ram[4424]  = 252;
  ram[4425]  = 250;
  ram[4426]  = 250;
  ram[4427]  = 253;
  ram[4428]  = 244;
  ram[4429]  = 242;
  ram[4430]  = 252;
  ram[4431]  = 250;
  ram[4432]  = 250;
  ram[4433]  = 250;
  ram[4434]  = 251;
  ram[4435]  = 252;
  ram[4436]  = 252;
  ram[4437]  = 253;
  ram[4438]  = 254;
  ram[4439]  = 243;
  ram[4440]  = 251;
  ram[4441]  = 252;
  ram[4442]  = 250;
  ram[4443]  = 250;
  ram[4444]  = 249;
  ram[4445]  = 248;
  ram[4446]  = 250;
  ram[4447]  = 250;
  ram[4448]  = 249;
  ram[4449]  = 247;
  ram[4450]  = 247;
  ram[4451]  = 131;
  ram[4452]  = 36;
  ram[4453]  = 3;
  ram[4454]  = 65;
  ram[4455]  = 232;
  ram[4456]  = 253;
  ram[4457]  = 252;
  ram[4458]  = 239;
  ram[4459]  = 253;
  ram[4460]  = 206;
  ram[4461]  = 0;
  ram[4462]  = 0;
  ram[4463]  = 0;
  ram[4464]  = 152;
  ram[4465]  = 255;
  ram[4466]  = 255;
  ram[4467]  = 255;
  ram[4468]  = 255;
  ram[4469]  = 255;
  ram[4470]  = 255;
  ram[4471]  = 255;
  ram[4472]  = 255;
  ram[4473]  = 255;
  ram[4474]  = 255;
  ram[4475]  = 255;
  ram[4476]  = 255;
  ram[4477]  = 255;
  ram[4478]  = 255;
  ram[4479]  = 255;
  ram[4480]  = 239;
  ram[4481]  = 245;
  ram[4482]  = 250;
  ram[4483]  = 251;
  ram[4484]  = 252;
  ram[4485]  = 251;
  ram[4486]  = 249;
  ram[4487]  = 251;
  ram[4488]  = 252;
  ram[4489]  = 252;
  ram[4490]  = 253;
  ram[4491]  = 255;
  ram[4492]  = 149;
  ram[4493]  = 0;
  ram[4494]  = 0;
  ram[4495]  = 20;
  ram[4496]  = 234;
  ram[4497]  = 254;
  ram[4498]  = 250;
  ram[4499]  = 250;
  ram[4500]  = 252;
  ram[4501]  = 255;
  ram[4502]  = 122;
  ram[4503]  = 13;
  ram[4504]  = 24;
  ram[4505]  = 54;
  ram[4506]  = 85;
  ram[4507]  = 104;
  ram[4508]  = 126;
  ram[4509]  = 179;
  ram[4510]  = 164;
  ram[4511]  = 0;
  ram[4512]  = 0;
  ram[4513]  = 0;
  ram[4514]  = 28;
  ram[4515]  = 234;
  ram[4516]  = 255;
  ram[4517]  = 252;
  ram[4518]  = 251;
  ram[4519]  = 252;
  ram[4520]  = 251;
  ram[4521]  = 252;
  ram[4522]  = 252;
  ram[4523]  = 253;
  ram[4524]  = 254;
  ram[4525]  = 247;
  ram[4526]  = 239;
  ram[4527]  = 251;
  ram[4528]  = 253;
  ram[4529]  = 253;
  ram[4530]  = 252;
  ram[4531]  = 252;
  ram[4532]  = 255;
  ram[4533]  = 186;
  ram[4534]  = 18;
  ram[4535]  = 0;
  ram[4536]  = 0;
  ram[4537]  = 0;
  ram[4538]  = 0;
  ram[4539]  = 0;
  ram[4540]  = 127;
  ram[4541]  = 255;
  ram[4542]  = 251;
  ram[4543]  = 250;
  ram[4544]  = 251;
  ram[4545]  = 249;
  ram[4546]  = 251;
  ram[4547]  = 253;
  ram[4548]  = 246;
  ram[4549]  = 244;
  ram[4550]  = 251;
  ram[4551]  = 249;
  ram[4552]  = 250;
  ram[4553]  = 251;
  ram[4554]  = 252;
  ram[4555]  = 252;
  ram[4556]  = 252;
  ram[4557]  = 253;
  ram[4558]  = 255;
  ram[4559]  = 242;
  ram[4560]  = 242;
  ram[4561]  = 240;
  ram[4562]  = 236;
  ram[4563]  = 239;
  ram[4564]  = 241;
  ram[4565]  = 239;
  ram[4566]  = 242;
  ram[4567]  = 240;
  ram[4568]  = 241;
  ram[4569]  = 231;
  ram[4570]  = 243;
  ram[4571]  = 255;
  ram[4572]  = 239;
  ram[4573]  = 206;
  ram[4574]  = 239;
  ram[4575]  = 251;
  ram[4576]  = 242;
  ram[4577]  = 242;
  ram[4578]  = 228;
  ram[4579]  = 235;
  ram[4580]  = 253;
  ram[4581]  = 93;
  ram[4582]  = 0;
  ram[4583]  = 13;
  ram[4584]  = 212;
  ram[4585]  = 248;
  ram[4586]  = 245;
  ram[4587]  = 242;
  ram[4588]  = 240;
  ram[4589]  = 230;
  ram[4590]  = 228;
  ram[4591]  = 238;
  ram[4592]  = 238;
  ram[4593]  = 238;
  ram[4594]  = 239;
  ram[4595]  = 238;
  ram[4596]  = 237;
  ram[4597]  = 238;
  ram[4598]  = 236;
  ram[4599]  = 236;
  ram[4600]  = 226;
  ram[4601]  = 232;
  ram[4602]  = 235;
  ram[4603]  = 239;
  ram[4604]  = 238;
  ram[4605]  = 237;
  ram[4606]  = 239;
  ram[4607]  = 243;
  ram[4608]  = 240;
  ram[4609]  = 240;
  ram[4610]  = 243;
  ram[4611]  = 238;
  ram[4612]  = 232;
  ram[4613]  = 86;
  ram[4614]  = 16;
  ram[4615]  = 120;
  ram[4616]  = 253;
  ram[4617]  = 242;
  ram[4618]  = 241;
  ram[4619]  = 237;
  ram[4620]  = 239;
  ram[4621]  = 247;
  ram[4622]  = 253;
  ram[4623]  = 208;
  ram[4624]  = 224;
  ram[4625]  = 248;
  ram[4626]  = 255;
  ram[4627]  = 255;
  ram[4628]  = 255;
  ram[4629]  = 255;
  ram[4630]  = 249;
  ram[4631]  = 71;
  ram[4632]  = 0;
  ram[4633]  = 0;
  ram[4634]  = 133;
  ram[4635]  = 251;
  ram[4636]  = 242;
  ram[4637]  = 242;
  ram[4638]  = 240;
  ram[4639]  = 240;
  ram[4640]  = 243;
  ram[4641]  = 241;
  ram[4642]  = 240;
  ram[4643]  = 244;
  ram[4644]  = 244;
  ram[4645]  = 233;
  ram[4646]  = 226;
  ram[4647]  = 241;
  ram[4648]  = 244;
  ram[4649]  = 244;
  ram[4650]  = 241;
  ram[4651]  = 240;
  ram[4652]  = 245;
  ram[4653]  = 254;
  ram[4654]  = 209;
  ram[4655]  = 109;
  ram[4656]  = 47;
  ram[4657]  = 7;
  ram[4658]  = 28;
  ram[4659]  = 127;
  ram[4660]  = 246;
  ram[4661]  = 244;
  ram[4662]  = 240;
  ram[4663]  = 238;
  ram[4664]  = 240;
  ram[4665]  = 240;
  ram[4666]  = 240;
  ram[4667]  = 241;
  ram[4668]  = 234;
  ram[4669]  = 231;
  ram[4670]  = 235;
  ram[4671]  = 234;
  ram[4672]  = 236;
  ram[4673]  = 240;
  ram[4674]  = 236;
  ram[4675]  = 240;
  ram[4676]  = 239;
  ram[4677]  = 239;
  ram[4678]  = 240;
  ram[4679]  = 231;
  ram[4680]  = 250;
  ram[4681]  = 251;
  ram[4682]  = 248;
  ram[4683]  = 249;
  ram[4684]  = 249;
  ram[4685]  = 249;
  ram[4686]  = 250;
  ram[4687]  = 251;
  ram[4688]  = 247;
  ram[4689]  = 236;
  ram[4690]  = 248;
  ram[4691]  = 253;
  ram[4692]  = 255;
  ram[4693]  = 255;
  ram[4694]  = 255;
  ram[4695]  = 251;
  ram[4696]  = 250;
  ram[4697]  = 250;
  ram[4698]  = 240;
  ram[4699]  = 243;
  ram[4700]  = 255;
  ram[4701]  = 247;
  ram[4702]  = 168;
  ram[4703]  = 174;
  ram[4704]  = 254;
  ram[4705]  = 249;
  ram[4706]  = 248;
  ram[4707]  = 248;
  ram[4708]  = 251;
  ram[4709]  = 240;
  ram[4710]  = 234;
  ram[4711]  = 246;
  ram[4712]  = 246;
  ram[4713]  = 246;
  ram[4714]  = 248;
  ram[4715]  = 242;
  ram[4716]  = 244;
  ram[4717]  = 246;
  ram[4718]  = 247;
  ram[4719]  = 249;
  ram[4720]  = 237;
  ram[4721]  = 242;
  ram[4722]  = 248;
  ram[4723]  = 249;
  ram[4724]  = 247;
  ram[4725]  = 246;
  ram[4726]  = 249;
  ram[4727]  = 250;
  ram[4728]  = 248;
  ram[4729]  = 248;
  ram[4730]  = 249;
  ram[4731]  = 241;
  ram[4732]  = 247;
  ram[4733]  = 255;
  ram[4734]  = 222;
  ram[4735]  = 255;
  ram[4736]  = 250;
  ram[4737]  = 249;
  ram[4738]  = 248;
  ram[4739]  = 245;
  ram[4740]  = 245;
  ram[4741]  = 250;
  ram[4742]  = 247;
  ram[4743]  = 248;
  ram[4744]  = 255;
  ram[4745]  = 250;
  ram[4746]  = 249;
  ram[4747]  = 250;
  ram[4748]  = 249;
  ram[4749]  = 248;
  ram[4750]  = 255;
  ram[4751]  = 229;
  ram[4752]  = 140;
  ram[4753]  = 196;
  ram[4754]  = 250;
  ram[4755]  = 241;
  ram[4756]  = 248;
  ram[4757]  = 249;
  ram[4758]  = 248;
  ram[4759]  = 246;
  ram[4760]  = 249;
  ram[4761]  = 247;
  ram[4762]  = 248;
  ram[4763]  = 249;
  ram[4764]  = 250;
  ram[4765]  = 242;
  ram[4766]  = 233;
  ram[4767]  = 248;
  ram[4768]  = 250;
  ram[4769]  = 248;
  ram[4770]  = 244;
  ram[4771]  = 247;
  ram[4772]  = 248;
  ram[4773]  = 245;
  ram[4774]  = 255;
  ram[4775]  = 255;
  ram[4776]  = 249;
  ram[4777]  = 215;
  ram[4778]  = 228;
  ram[4779]  = 255;
  ram[4780]  = 249;
  ram[4781]  = 245;
  ram[4782]  = 246;
  ram[4783]  = 245;
  ram[4784]  = 246;
  ram[4785]  = 248;
  ram[4786]  = 248;
  ram[4787]  = 248;
  ram[4788]  = 240;
  ram[4789]  = 236;
  ram[4790]  = 246;
  ram[4791]  = 243;
  ram[4792]  = 243;
  ram[4793]  = 246;
  ram[4794]  = 244;
  ram[4795]  = 244;
  ram[4796]  = 245;
  ram[4797]  = 246;
  ram[4798]  = 246;
  ram[4799]  = 237;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
