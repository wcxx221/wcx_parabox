module rom_tui1(clock, address, q);     // ROM-stored RGB bitmap for display region 1
input clock;
output [7:0] q;
input [12:0] address;
reg [7:0] dout;
reg [7:0] ram [8191:0];
assign q = dout;

initial begin
  ram[0]  = 255;
  ram[1]  = 255;
  ram[2]  = 255;
  ram[3]  = 255;
  ram[4]  = 255;
  ram[5]  = 255;
  ram[6]  = 255;
  ram[7]  = 255;
  ram[8]  = 255;
  ram[9]  = 255;
  ram[10]  = 255;
  ram[11]  = 255;
  ram[12]  = 255;
  ram[13]  = 255;
  ram[14]  = 255;
  ram[15]  = 255;
  ram[16]  = 255;
  ram[17]  = 255;
  ram[18]  = 255;
  ram[19]  = 255;
  ram[20]  = 255;
  ram[21]  = 255;
  ram[22]  = 255;
  ram[23]  = 255;
  ram[24]  = 255;
  ram[25]  = 255;
  ram[26]  = 255;
  ram[27]  = 255;
  ram[28]  = 255;
  ram[29]  = 255;
  ram[30]  = 255;
  ram[31]  = 255;
  ram[32]  = 255;
  ram[33]  = 255;
  ram[34]  = 255;
  ram[35]  = 255;
  ram[36]  = 255;
  ram[37]  = 255;
  ram[38]  = 255;
  ram[39]  = 255;
  ram[40]  = 255;
  ram[41]  = 255;
  ram[42]  = 255;
  ram[43]  = 255;
  ram[44]  = 255;
  ram[45]  = 255;
  ram[46]  = 255;
  ram[47]  = 255;
  ram[48]  = 255;
  ram[49]  = 255;
  ram[50]  = 255;
  ram[51]  = 255;
  ram[52]  = 255;
  ram[53]  = 255;
  ram[54]  = 255;
  ram[55]  = 255;
  ram[56]  = 255;
  ram[57]  = 255;
  ram[58]  = 255;
  ram[59]  = 255;
  ram[60]  = 255;
  ram[61]  = 255;
  ram[62]  = 255;
  ram[63]  = 255;
  ram[64]  = 255;
  ram[65]  = 255;
  ram[66]  = 255;
  ram[67]  = 255;
  ram[68]  = 255;
  ram[69]  = 255;
  ram[70]  = 255;
  ram[71]  = 255;
  ram[72]  = 255;
  ram[73]  = 255;
  ram[74]  = 255;
  ram[75]  = 255;
  ram[76]  = 255;
  ram[77]  = 255;
  ram[78]  = 255;
  ram[79]  = 255;
  ram[80]  = 255;
  ram[81]  = 255;
  ram[82]  = 255;
  ram[83]  = 255;
  ram[84]  = 255;
  ram[85]  = 255;
  ram[86]  = 255;
  ram[87]  = 255;
  ram[88]  = 255;
  ram[89]  = 255;
  ram[90]  = 255;
  ram[91]  = 255;
  ram[92]  = 255;
  ram[93]  = 255;
  ram[94]  = 255;
  ram[95]  = 255;
  ram[96]  = 255;
  ram[97]  = 255;
  ram[98]  = 255;
  ram[99]  = 255;
  ram[100]  = 255;
  ram[101]  = 255;
  ram[102]  = 255;
  ram[103]  = 255;
  ram[104]  = 255;
  ram[105]  = 255;
  ram[106]  = 255;
  ram[107]  = 255;
  ram[108]  = 255;
  ram[109]  = 255;
  ram[110]  = 255;
  ram[111]  = 255;
  ram[112]  = 255;
  ram[113]  = 255;
  ram[114]  = 255;
  ram[115]  = 255;
  ram[116]  = 255;
  ram[117]  = 255;
  ram[118]  = 255;
  ram[119]  = 255;
  ram[120]  = 255;
  ram[121]  = 255;
  ram[122]  = 255;
  ram[123]  = 255;
  ram[124]  = 255;
  ram[125]  = 255;
  ram[126]  = 255;
  ram[127]  = 255;
  ram[128]  = 255;
  ram[129]  = 255;
  ram[130]  = 255;
  ram[131]  = 255;
  ram[132]  = 255;
  ram[133]  = 255;
  ram[134]  = 255;
  ram[135]  = 255;
  ram[136]  = 255;
  ram[137]  = 255;
  ram[138]  = 255;
  ram[139]  = 255;
  ram[140]  = 255;
  ram[141]  = 255;
  ram[142]  = 255;
  ram[143]  = 255;
  ram[144]  = 255;
  ram[145]  = 255;
  ram[146]  = 255;
  ram[147]  = 255;
  ram[148]  = 255;
  ram[149]  = 255;
  ram[150]  = 255;
  ram[151]  = 255;
  ram[152]  = 255;
  ram[153]  = 255;
  ram[154]  = 255;
  ram[155]  = 255;
  ram[156]  = 255;
  ram[157]  = 255;
  ram[158]  = 255;
  ram[159]  = 255;
  ram[160]  = 255;
  ram[161]  = 255;
  ram[162]  = 255;
  ram[163]  = 255;
  ram[164]  = 255;
  ram[165]  = 255;
  ram[166]  = 255;
  ram[167]  = 255;
  ram[168]  = 255;
  ram[169]  = 255;
  ram[170]  = 255;
  ram[171]  = 255;
  ram[172]  = 255;
  ram[173]  = 255;
  ram[174]  = 255;
  ram[175]  = 255;
  ram[176]  = 255;
  ram[177]  = 255;
  ram[178]  = 255;
  ram[179]  = 255;
  ram[180]  = 255;
  ram[181]  = 255;
  ram[182]  = 255;
  ram[183]  = 255;
  ram[184]  = 255;
  ram[185]  = 255;
  ram[186]  = 255;
  ram[187]  = 255;
  ram[188]  = 255;
  ram[189]  = 255;
  ram[190]  = 255;
  ram[191]  = 255;
  ram[192]  = 255;
  ram[193]  = 255;
  ram[194]  = 255;
  ram[195]  = 255;
  ram[196]  = 255;
  ram[197]  = 255;
  ram[198]  = 255;
  ram[199]  = 255;
  ram[200]  = 255;
  ram[201]  = 255;
  ram[202]  = 255;
  ram[203]  = 255;
  ram[204]  = 255;
  ram[205]  = 255;
  ram[206]  = 255;
  ram[207]  = 255;
  ram[208]  = 255;
  ram[209]  = 255;
  ram[210]  = 255;
  ram[211]  = 255;
  ram[212]  = 255;
  ram[213]  = 255;
  ram[214]  = 255;
  ram[215]  = 255;
  ram[216]  = 255;
  ram[217]  = 255;
  ram[218]  = 255;
  ram[219]  = 255;
  ram[220]  = 255;
  ram[221]  = 255;
  ram[222]  = 255;
  ram[223]  = 255;
  ram[224]  = 255;
  ram[225]  = 255;
  ram[226]  = 255;
  ram[227]  = 255;
  ram[228]  = 255;
  ram[229]  = 255;
  ram[230]  = 255;
  ram[231]  = 255;
  ram[232]  = 255;
  ram[233]  = 255;
  ram[234]  = 255;
  ram[235]  = 255;
  ram[236]  = 255;
  ram[237]  = 255;
  ram[238]  = 255;
  ram[239]  = 255;
  ram[240]  = 255;
  ram[241]  = 255;
  ram[242]  = 255;
  ram[243]  = 255;
  ram[244]  = 255;
  ram[245]  = 255;
  ram[246]  = 255;
  ram[247]  = 255;
  ram[248]  = 255;
  ram[249]  = 255;
  ram[250]  = 255;
  ram[251]  = 255;
  ram[252]  = 255;
  ram[253]  = 255;
  ram[254]  = 255;
  ram[255]  = 255;
  ram[256]  = 255;
  ram[257]  = 255;
  ram[258]  = 255;
  ram[259]  = 255;
  ram[260]  = 255;
  ram[261]  = 255;
  ram[262]  = 255;
  ram[263]  = 255;
  ram[264]  = 255;
  ram[265]  = 255;
  ram[266]  = 255;
  ram[267]  = 255;
  ram[268]  = 255;
  ram[269]  = 255;
  ram[270]  = 255;
  ram[271]  = 255;
  ram[272]  = 255;
  ram[273]  = 255;
  ram[274]  = 255;
  ram[275]  = 255;
  ram[276]  = 255;
  ram[277]  = 255;
  ram[278]  = 255;
  ram[279]  = 255;
  ram[280]  = 255;
  ram[281]  = 255;
  ram[282]  = 255;
  ram[283]  = 255;
  ram[284]  = 255;
  ram[285]  = 255;
  ram[286]  = 255;
  ram[287]  = 255;
  ram[288]  = 255;
  ram[289]  = 255;
  ram[290]  = 255;
  ram[291]  = 255;
  ram[292]  = 255;
  ram[293]  = 255;
  ram[294]  = 255;
  ram[295]  = 255;
  ram[296]  = 255;
  ram[297]  = 255;
  ram[298]  = 255;
  ram[299]  = 255;
  ram[300]  = 255;
  ram[301]  = 255;
  ram[302]  = 255;
  ram[303]  = 255;
  ram[304]  = 255;
  ram[305]  = 255;
  ram[306]  = 255;
  ram[307]  = 255;
  ram[308]  = 255;
  ram[309]  = 255;
  ram[310]  = 255;
  ram[311]  = 255;
  ram[312]  = 255;
  ram[313]  = 255;
  ram[314]  = 255;
  ram[315]  = 255;
  ram[316]  = 255;
  ram[317]  = 255;
  ram[318]  = 255;
  ram[319]  = 255;
  ram[320]  = 255;
  ram[321]  = 255;
  ram[322]  = 255;
  ram[323]  = 255;
  ram[324]  = 255;
  ram[325]  = 255;
  ram[326]  = 255;
  ram[327]  = 255;
  ram[328]  = 255;
  ram[329]  = 255;
  ram[330]  = 255;
  ram[331]  = 255;
  ram[332]  = 255;
  ram[333]  = 255;
  ram[334]  = 255;
  ram[335]  = 255;
  ram[336]  = 255;
  ram[337]  = 255;
  ram[338]  = 255;
  ram[339]  = 255;
  ram[340]  = 255;
  ram[341]  = 255;
  ram[342]  = 255;
  ram[343]  = 255;
  ram[344]  = 255;
  ram[345]  = 255;
  ram[346]  = 255;
  ram[347]  = 255;
  ram[348]  = 255;
  ram[349]  = 255;
  ram[350]  = 255;
  ram[351]  = 255;
  ram[352]  = 255;
  ram[353]  = 255;
  ram[354]  = 255;
  ram[355]  = 255;
  ram[356]  = 255;
  ram[357]  = 255;
  ram[358]  = 255;
  ram[359]  = 255;
  ram[360]  = 255;
  ram[361]  = 255;
  ram[362]  = 255;
  ram[363]  = 255;
  ram[364]  = 255;
  ram[365]  = 255;
  ram[366]  = 255;
  ram[367]  = 255;
  ram[368]  = 255;
  ram[369]  = 255;
  ram[370]  = 255;
  ram[371]  = 255;
  ram[372]  = 255;
  ram[373]  = 255;
  ram[374]  = 255;
  ram[375]  = 255;
  ram[376]  = 255;
  ram[377]  = 255;
  ram[378]  = 255;
  ram[379]  = 255;
  ram[380]  = 255;
  ram[381]  = 255;
  ram[382]  = 255;
  ram[383]  = 255;
  ram[384]  = 255;
  ram[385]  = 255;
  ram[386]  = 255;
  ram[387]  = 255;
  ram[388]  = 255;
  ram[389]  = 255;
  ram[390]  = 255;
  ram[391]  = 255;
  ram[392]  = 255;
  ram[393]  = 255;
  ram[394]  = 255;
  ram[395]  = 255;
  ram[396]  = 255;
  ram[397]  = 255;
  ram[398]  = 255;
  ram[399]  = 255;
  ram[400]  = 255;
  ram[401]  = 255;
  ram[402]  = 255;
  ram[403]  = 255;
  ram[404]  = 255;
  ram[405]  = 255;
  ram[406]  = 255;
  ram[407]  = 255;
  ram[408]  = 255;
  ram[409]  = 255;
  ram[410]  = 255;
  ram[411]  = 255;
  ram[412]  = 255;
  ram[413]  = 255;
  ram[414]  = 255;
  ram[415]  = 255;
  ram[416]  = 255;
  ram[417]  = 255;
  ram[418]  = 255;
  ram[419]  = 255;
  ram[420]  = 255;
  ram[421]  = 255;
  ram[422]  = 255;
  ram[423]  = 255;
  ram[424]  = 255;
  ram[425]  = 255;
  ram[426]  = 255;
  ram[427]  = 255;
  ram[428]  = 255;
  ram[429]  = 255;
  ram[430]  = 255;
  ram[431]  = 255;
  ram[432]  = 255;
  ram[433]  = 255;
  ram[434]  = 255;
  ram[435]  = 255;
  ram[436]  = 255;
  ram[437]  = 255;
  ram[438]  = 255;
  ram[439]  = 255;
  ram[440]  = 255;
  ram[441]  = 255;
  ram[442]  = 255;
  ram[443]  = 255;
  ram[444]  = 255;
  ram[445]  = 255;
  ram[446]  = 255;
  ram[447]  = 255;
  ram[448]  = 255;
  ram[449]  = 255;
  ram[450]  = 255;
  ram[451]  = 255;
  ram[452]  = 255;
  ram[453]  = 255;
  ram[454]  = 255;
  ram[455]  = 255;
  ram[456]  = 255;
  ram[457]  = 255;
  ram[458]  = 255;
  ram[459]  = 255;
  ram[460]  = 255;
  ram[461]  = 255;
  ram[462]  = 255;
  ram[463]  = 255;
  ram[464]  = 255;
  ram[465]  = 255;
  ram[466]  = 255;
  ram[467]  = 255;
  ram[468]  = 255;
  ram[469]  = 255;
  ram[470]  = 255;
  ram[471]  = 255;
  ram[472]  = 255;
  ram[473]  = 255;
  ram[474]  = 255;
  ram[475]  = 255;
  ram[476]  = 255;
  ram[477]  = 255;
  ram[478]  = 255;
  ram[479]  = 255;
  ram[480]  = 255;
  ram[481]  = 255;
  ram[482]  = 255;
  ram[483]  = 255;
  ram[484]  = 255;
  ram[485]  = 255;
  ram[486]  = 255;
  ram[487]  = 255;
  ram[488]  = 255;
  ram[489]  = 255;
  ram[490]  = 255;
  ram[491]  = 255;
  ram[492]  = 255;
  ram[493]  = 255;
  ram[494]  = 255;
  ram[495]  = 255;
  ram[496]  = 255;
  ram[497]  = 255;
  ram[498]  = 255;
  ram[499]  = 255;
  ram[500]  = 255;
  ram[501]  = 255;
  ram[502]  = 255;
  ram[503]  = 255;
  ram[504]  = 255;
  ram[505]  = 255;
  ram[506]  = 255;
  ram[507]  = 255;
  ram[508]  = 255;
  ram[509]  = 255;
  ram[510]  = 255;
  ram[511]  = 255;
  ram[512]  = 255;
  ram[513]  = 255;
  ram[514]  = 255;
  ram[515]  = 255;
  ram[516]  = 255;
  ram[517]  = 255;
  ram[518]  = 255;
  ram[519]  = 255;
  ram[520]  = 255;
  ram[521]  = 255;
  ram[522]  = 255;
  ram[523]  = 255;
  ram[524]  = 255;
  ram[525]  = 255;
  ram[526]  = 255;
  ram[527]  = 255;
  ram[528]  = 255;
  ram[529]  = 255;
  ram[530]  = 255;
  ram[531]  = 255;
  ram[532]  = 255;
  ram[533]  = 255;
  ram[534]  = 255;
  ram[535]  = 255;
  ram[536]  = 255;
  ram[537]  = 255;
  ram[538]  = 255;
  ram[539]  = 255;
  ram[540]  = 255;
  ram[541]  = 255;
  ram[542]  = 255;
  ram[543]  = 255;
  ram[544]  = 255;
  ram[545]  = 255;
  ram[546]  = 255;
  ram[547]  = 255;
  ram[548]  = 255;
  ram[549]  = 255;
  ram[550]  = 255;
  ram[551]  = 255;
  ram[552]  = 255;
  ram[553]  = 255;
  ram[554]  = 255;
  ram[555]  = 255;
  ram[556]  = 255;
  ram[557]  = 255;
  ram[558]  = 255;
  ram[559]  = 255;
  ram[560]  = 255;
  ram[561]  = 255;
  ram[562]  = 255;
  ram[563]  = 255;
  ram[564]  = 255;
  ram[565]  = 255;
  ram[566]  = 255;
  ram[567]  = 255;
  ram[568]  = 255;
  ram[569]  = 255;
  ram[570]  = 255;
  ram[571]  = 255;
  ram[572]  = 255;
  ram[573]  = 255;
  ram[574]  = 255;
  ram[575]  = 255;
  ram[576]  = 255;
  ram[577]  = 255;
  ram[578]  = 255;
  ram[579]  = 255;
  ram[580]  = 255;
  ram[581]  = 255;
  ram[582]  = 255;
  ram[583]  = 255;
  ram[584]  = 255;
  ram[585]  = 255;
  ram[586]  = 255;
  ram[587]  = 255;
  ram[588]  = 255;
  ram[589]  = 255;
  ram[590]  = 255;
  ram[591]  = 255;
  ram[592]  = 255;
  ram[593]  = 255;
  ram[594]  = 255;
  ram[595]  = 255;
  ram[596]  = 255;
  ram[597]  = 255;
  ram[598]  = 255;
  ram[599]  = 255;
  ram[600]  = 255;
  ram[601]  = 255;
  ram[602]  = 255;
  ram[603]  = 255;
  ram[604]  = 255;
  ram[605]  = 255;
  ram[606]  = 255;
  ram[607]  = 255;
  ram[608]  = 255;
  ram[609]  = 255;
  ram[610]  = 255;
  ram[611]  = 255;
  ram[612]  = 255;
  ram[613]  = 255;
  ram[614]  = 255;
  ram[615]  = 255;
  ram[616]  = 255;
  ram[617]  = 255;
  ram[618]  = 255;
  ram[619]  = 255;
  ram[620]  = 255;
  ram[621]  = 255;
  ram[622]  = 255;
  ram[623]  = 255;
  ram[624]  = 255;
  ram[625]  = 255;
  ram[626]  = 255;
  ram[627]  = 255;
  ram[628]  = 255;
  ram[629]  = 255;
  ram[630]  = 255;
  ram[631]  = 255;
  ram[632]  = 255;
  ram[633]  = 255;
  ram[634]  = 255;
  ram[635]  = 255;
  ram[636]  = 255;
  ram[637]  = 255;
  ram[638]  = 255;
  ram[639]  = 255;
  ram[640]  = 255;
  ram[641]  = 255;
  ram[642]  = 255;
  ram[643]  = 255;
  ram[644]  = 255;
  ram[645]  = 255;
  ram[646]  = 255;
  ram[647]  = 255;
  ram[648]  = 255;
  ram[649]  = 255;
  ram[650]  = 255;
  ram[651]  = 255;
  ram[652]  = 255;
  ram[653]  = 255;
  ram[654]  = 255;
  ram[655]  = 255;
  ram[656]  = 255;
  ram[657]  = 255;
  ram[658]  = 255;
  ram[659]  = 255;
  ram[660]  = 255;
  ram[661]  = 255;
  ram[662]  = 255;
  ram[663]  = 255;
  ram[664]  = 255;
  ram[665]  = 255;
  ram[666]  = 255;
  ram[667]  = 255;
  ram[668]  = 255;
  ram[669]  = 255;
  ram[670]  = 255;
  ram[671]  = 255;
  ram[672]  = 255;
  ram[673]  = 255;
  ram[674]  = 255;
  ram[675]  = 255;
  ram[676]  = 255;
  ram[677]  = 255;
  ram[678]  = 255;
  ram[679]  = 255;
  ram[680]  = 255;
  ram[681]  = 255;
  ram[682]  = 255;
  ram[683]  = 255;
  ram[684]  = 255;
  ram[685]  = 255;
  ram[686]  = 255;
  ram[687]  = 255;
  ram[688]  = 255;
  ram[689]  = 255;
  ram[690]  = 255;
  ram[691]  = 255;
  ram[692]  = 255;
  ram[693]  = 255;
  ram[694]  = 255;
  ram[695]  = 255;
  ram[696]  = 255;
  ram[697]  = 255;
  ram[698]  = 255;
  ram[699]  = 255;
  ram[700]  = 255;
  ram[701]  = 255;
  ram[702]  = 255;
  ram[703]  = 255;
  ram[704]  = 255;
  ram[705]  = 255;
  ram[706]  = 255;
  ram[707]  = 255;
  ram[708]  = 255;
  ram[709]  = 255;
  ram[710]  = 255;
  ram[711]  = 255;
  ram[712]  = 255;
  ram[713]  = 255;
  ram[714]  = 255;
  ram[715]  = 255;
  ram[716]  = 255;
  ram[717]  = 255;
  ram[718]  = 255;
  ram[719]  = 255;
  ram[720]  = 255;
  ram[721]  = 255;
  ram[722]  = 255;
  ram[723]  = 255;
  ram[724]  = 255;
  ram[725]  = 255;
  ram[726]  = 255;
  ram[727]  = 255;
  ram[728]  = 255;
  ram[729]  = 255;
  ram[730]  = 255;
  ram[731]  = 255;
  ram[732]  = 255;
  ram[733]  = 255;
  ram[734]  = 255;
  ram[735]  = 255;
  ram[736]  = 255;
  ram[737]  = 255;
  ram[738]  = 255;
  ram[739]  = 255;
  ram[740]  = 255;
  ram[741]  = 255;
  ram[742]  = 255;
  ram[743]  = 255;
  ram[744]  = 255;
  ram[745]  = 255;
  ram[746]  = 255;
  ram[747]  = 255;
  ram[748]  = 255;
  ram[749]  = 255;
  ram[750]  = 255;
  ram[751]  = 255;
  ram[752]  = 255;
  ram[753]  = 255;
  ram[754]  = 255;
  ram[755]  = 255;
  ram[756]  = 255;
  ram[757]  = 255;
  ram[758]  = 255;
  ram[759]  = 255;
  ram[760]  = 255;
  ram[761]  = 255;
  ram[762]  = 255;
  ram[763]  = 255;
  ram[764]  = 255;
  ram[765]  = 255;
  ram[766]  = 255;
  ram[767]  = 255;
  ram[768]  = 255;
  ram[769]  = 255;
  ram[770]  = 255;
  ram[771]  = 255;
  ram[772]  = 255;
  ram[773]  = 255;
  ram[774]  = 255;
  ram[775]  = 255;
  ram[776]  = 255;
  ram[777]  = 255;
  ram[778]  = 255;
  ram[779]  = 255;
  ram[780]  = 255;
  ram[781]  = 255;
  ram[782]  = 255;
  ram[783]  = 255;
  ram[784]  = 255;
  ram[785]  = 255;
  ram[786]  = 255;
  ram[787]  = 255;
  ram[788]  = 255;
  ram[789]  = 255;
  ram[790]  = 255;
  ram[791]  = 255;
  ram[792]  = 255;
  ram[793]  = 255;
  ram[794]  = 255;
  ram[795]  = 255;
  ram[796]  = 255;
  ram[797]  = 255;
  ram[798]  = 255;
  ram[799]  = 255;
  ram[800]  = 255;
  ram[801]  = 255;
  ram[802]  = 255;
  ram[803]  = 255;
  ram[804]  = 255;
  ram[805]  = 255;
  ram[806]  = 255;
  ram[807]  = 255;
  ram[808]  = 255;
  ram[809]  = 255;
  ram[810]  = 255;
  ram[811]  = 255;
  ram[812]  = 255;
  ram[813]  = 255;
  ram[814]  = 255;
  ram[815]  = 255;
  ram[816]  = 255;
  ram[817]  = 255;
  ram[818]  = 255;
  ram[819]  = 255;
  ram[820]  = 255;
  ram[821]  = 255;
  ram[822]  = 255;
  ram[823]  = 255;
  ram[824]  = 255;
  ram[825]  = 255;
  ram[826]  = 255;
  ram[827]  = 255;
  ram[828]  = 255;
  ram[829]  = 255;
  ram[830]  = 255;
  ram[831]  = 255;
  ram[832]  = 255;
  ram[833]  = 255;
  ram[834]  = 255;
  ram[835]  = 255;
  ram[836]  = 255;
  ram[837]  = 255;
  ram[838]  = 255;
  ram[839]  = 255;
  ram[840]  = 255;
  ram[841]  = 255;
  ram[842]  = 255;
  ram[843]  = 255;
  ram[844]  = 255;
  ram[845]  = 255;
  ram[846]  = 255;
  ram[847]  = 255;
  ram[848]  = 255;
  ram[849]  = 255;
  ram[850]  = 255;
  ram[851]  = 255;
  ram[852]  = 255;
  ram[853]  = 255;
  ram[854]  = 255;
  ram[855]  = 255;
  ram[856]  = 255;
  ram[857]  = 255;
  ram[858]  = 255;
  ram[859]  = 255;
  ram[860]  = 255;
  ram[861]  = 255;
  ram[862]  = 255;
  ram[863]  = 255;
  ram[864]  = 255;
  ram[865]  = 255;
  ram[866]  = 255;
  ram[867]  = 255;
  ram[868]  = 255;
  ram[869]  = 255;
  ram[870]  = 255;
  ram[871]  = 255;
  ram[872]  = 255;
  ram[873]  = 255;
  ram[874]  = 255;
  ram[875]  = 255;
  ram[876]  = 255;
  ram[877]  = 255;
  ram[878]  = 255;
  ram[879]  = 255;
  ram[880]  = 255;
  ram[881]  = 255;
  ram[882]  = 255;
  ram[883]  = 255;
  ram[884]  = 255;
  ram[885]  = 255;
  ram[886]  = 255;
  ram[887]  = 255;
  ram[888]  = 255;
  ram[889]  = 255;
  ram[890]  = 255;
  ram[891]  = 255;
  ram[892]  = 255;
  ram[893]  = 255;
  ram[894]  = 255;
  ram[895]  = 255;
  ram[896]  = 255;
  ram[897]  = 255;
  ram[898]  = 255;
  ram[899]  = 255;
  ram[900]  = 255;
  ram[901]  = 255;
  ram[902]  = 255;
  ram[903]  = 255;
  ram[904]  = 255;
  ram[905]  = 255;
  ram[906]  = 255;
  ram[907]  = 255;
  ram[908]  = 255;
  ram[909]  = 255;
  ram[910]  = 255;
  ram[911]  = 255;
  ram[912]  = 255;
  ram[913]  = 255;
  ram[914]  = 255;
  ram[915]  = 221;
  ram[916]  = 195;
  ram[917]  = 255;
  ram[918]  = 255;
  ram[919]  = 255;
  ram[920]  = 255;
  ram[921]  = 255;
  ram[922]  = 255;
  ram[923]  = 255;
  ram[924]  = 255;
  ram[925]  = 255;
  ram[926]  = 255;
  ram[927]  = 221;
  ram[928]  = 181;
  ram[929]  = 255;
  ram[930]  = 255;
  ram[931]  = 255;
  ram[932]  = 255;
  ram[933]  = 255;
  ram[934]  = 255;
  ram[935]  = 255;
  ram[936]  = 255;
  ram[937]  = 255;
  ram[938]  = 255;
  ram[939]  = 255;
  ram[940]  = 255;
  ram[941]  = 255;
  ram[942]  = 255;
  ram[943]  = 255;
  ram[944]  = 255;
  ram[945]  = 255;
  ram[946]  = 255;
  ram[947]  = 255;
  ram[948]  = 255;
  ram[949]  = 255;
  ram[950]  = 255;
  ram[951]  = 255;
  ram[952]  = 255;
  ram[953]  = 255;
  ram[954]  = 255;
  ram[955]  = 255;
  ram[956]  = 255;
  ram[957]  = 255;
  ram[958]  = 255;
  ram[959]  = 255;
  ram[960]  = 255;
  ram[961]  = 255;
  ram[962]  = 255;
  ram[963]  = 255;
  ram[964]  = 255;
  ram[965]  = 255;
  ram[966]  = 255;
  ram[967]  = 255;
  ram[968]  = 255;
  ram[969]  = 255;
  ram[970]  = 255;
  ram[971]  = 255;
  ram[972]  = 255;
  ram[973]  = 255;
  ram[974]  = 255;
  ram[975]  = 255;
  ram[976]  = 255;
  ram[977]  = 255;
  ram[978]  = 255;
  ram[979]  = 255;
  ram[980]  = 255;
  ram[981]  = 255;
  ram[982]  = 255;
  ram[983]  = 255;
  ram[984]  = 255;
  ram[985]  = 255;
  ram[986]  = 255;
  ram[987]  = 255;
  ram[988]  = 255;
  ram[989]  = 255;
  ram[990]  = 255;
  ram[991]  = 255;
  ram[992]  = 255;
  ram[993]  = 255;
  ram[994]  = 255;
  ram[995]  = 255;
  ram[996]  = 255;
  ram[997]  = 255;
  ram[998]  = 255;
  ram[999]  = 255;
  ram[1000]  = 255;
  ram[1001]  = 255;
  ram[1002]  = 255;
  ram[1003]  = 255;
  ram[1004]  = 255;
  ram[1005]  = 255;
  ram[1006]  = 255;
  ram[1007]  = 255;
  ram[1008]  = 255;
  ram[1009]  = 255;
  ram[1010]  = 255;
  ram[1011]  = 255;
  ram[1012]  = 255;
  ram[1013]  = 255;
  ram[1014]  = 255;
  ram[1015]  = 255;
  ram[1016]  = 255;
  ram[1017]  = 255;
  ram[1018]  = 255;
  ram[1019]  = 255;
  ram[1020]  = 255;
  ram[1021]  = 255;
  ram[1022]  = 255;
  ram[1023]  = 255;
  ram[1024]  = 255;
  ram[1025]  = 255;
  ram[1026]  = 255;
  ram[1027]  = 255;
  ram[1028]  = 255;
  ram[1029]  = 255;
  ram[1030]  = 255;
  ram[1031]  = 255;
  ram[1032]  = 255;
  ram[1033]  = 255;
  ram[1034]  = 255;
  ram[1035]  = 137;
  ram[1036]  = 0;
  ram[1037]  = 105;
  ram[1038]  = 255;
  ram[1039]  = 255;
  ram[1040]  = 255;
  ram[1041]  = 255;
  ram[1042]  = 255;
  ram[1043]  = 255;
  ram[1044]  = 255;
  ram[1045]  = 255;
  ram[1046]  = 255;
  ram[1047]  = 105;
  ram[1048]  = 0;
  ram[1049]  = 52;
  ram[1050]  = 255;
  ram[1051]  = 255;
  ram[1052]  = 255;
  ram[1053]  = 255;
  ram[1054]  = 255;
  ram[1055]  = 255;
  ram[1056]  = 255;
  ram[1057]  = 255;
  ram[1058]  = 255;
  ram[1059]  = 255;
  ram[1060]  = 255;
  ram[1061]  = 255;
  ram[1062]  = 255;
  ram[1063]  = 255;
  ram[1064]  = 255;
  ram[1065]  = 255;
  ram[1066]  = 255;
  ram[1067]  = 255;
  ram[1068]  = 255;
  ram[1069]  = 255;
  ram[1070]  = 255;
  ram[1071]  = 255;
  ram[1072]  = 255;
  ram[1073]  = 255;
  ram[1074]  = 255;
  ram[1075]  = 255;
  ram[1076]  = 255;
  ram[1077]  = 255;
  ram[1078]  = 255;
  ram[1079]  = 255;
  ram[1080]  = 255;
  ram[1081]  = 255;
  ram[1082]  = 255;
  ram[1083]  = 255;
  ram[1084]  = 255;
  ram[1085]  = 255;
  ram[1086]  = 255;
  ram[1087]  = 255;
  ram[1088]  = 255;
  ram[1089]  = 255;
  ram[1090]  = 255;
  ram[1091]  = 181;
  ram[1092]  = 122;
  ram[1093]  = 71;
  ram[1094]  = 71;
  ram[1095]  = 71;
  ram[1096]  = 71;
  ram[1097]  = 137;
  ram[1098]  = 181;
  ram[1099]  = 236;
  ram[1100]  = 255;
  ram[1101]  = 255;
  ram[1102]  = 255;
  ram[1103]  = 255;
  ram[1104]  = 255;
  ram[1105]  = 255;
  ram[1106]  = 255;
  ram[1107]  = 255;
  ram[1108]  = 255;
  ram[1109]  = 255;
  ram[1110]  = 255;
  ram[1111]  = 255;
  ram[1112]  = 255;
  ram[1113]  = 255;
  ram[1114]  = 255;
  ram[1115]  = 255;
  ram[1116]  = 255;
  ram[1117]  = 255;
  ram[1118]  = 167;
  ram[1119]  = 137;
  ram[1120]  = 137;
  ram[1121]  = 137;
  ram[1122]  = 137;
  ram[1123]  = 137;
  ram[1124]  = 137;
  ram[1125]  = 137;
  ram[1126]  = 137;
  ram[1127]  = 137;
  ram[1128]  = 137;
  ram[1129]  = 137;
  ram[1130]  = 137;
  ram[1131]  = 137;
  ram[1132]  = 137;
  ram[1133]  = 137;
  ram[1134]  = 137;
  ram[1135]  = 137;
  ram[1136]  = 137;
  ram[1137]  = 137;
  ram[1138]  = 137;
  ram[1139]  = 137;
  ram[1140]  = 137;
  ram[1141]  = 167;
  ram[1142]  = 255;
  ram[1143]  = 255;
  ram[1144]  = 255;
  ram[1145]  = 255;
  ram[1146]  = 255;
  ram[1147]  = 255;
  ram[1148]  = 255;
  ram[1149]  = 255;
  ram[1150]  = 255;
  ram[1151]  = 255;
  ram[1152]  = 255;
  ram[1153]  = 255;
  ram[1154]  = 255;
  ram[1155]  = 87;
  ram[1156]  = 0;
  ram[1157]  = 137;
  ram[1158]  = 255;
  ram[1159]  = 255;
  ram[1160]  = 255;
  ram[1161]  = 255;
  ram[1162]  = 255;
  ram[1163]  = 255;
  ram[1164]  = 255;
  ram[1165]  = 255;
  ram[1166]  = 221;
  ram[1167]  = 0;
  ram[1168]  = 0;
  ram[1169]  = 167;
  ram[1170]  = 255;
  ram[1171]  = 255;
  ram[1172]  = 255;
  ram[1173]  = 255;
  ram[1174]  = 255;
  ram[1175]  = 255;
  ram[1176]  = 255;
  ram[1177]  = 255;
  ram[1178]  = 255;
  ram[1179]  = 255;
  ram[1180]  = 255;
  ram[1181]  = 255;
  ram[1182]  = 255;
  ram[1183]  = 255;
  ram[1184]  = 255;
  ram[1185]  = 255;
  ram[1186]  = 255;
  ram[1187]  = 255;
  ram[1188]  = 255;
  ram[1189]  = 255;
  ram[1190]  = 255;
  ram[1191]  = 255;
  ram[1192]  = 255;
  ram[1193]  = 255;
  ram[1194]  = 255;
  ram[1195]  = 255;
  ram[1196]  = 255;
  ram[1197]  = 255;
  ram[1198]  = 255;
  ram[1199]  = 255;
  ram[1200]  = 255;
  ram[1201]  = 255;
  ram[1202]  = 255;
  ram[1203]  = 255;
  ram[1204]  = 255;
  ram[1205]  = 255;
  ram[1206]  = 255;
  ram[1207]  = 255;
  ram[1208]  = 255;
  ram[1209]  = 137;
  ram[1210]  = 17;
  ram[1211]  = 0;
  ram[1212]  = 0;
  ram[1213]  = 0;
  ram[1214]  = 0;
  ram[1215]  = 0;
  ram[1216]  = 0;
  ram[1217]  = 0;
  ram[1218]  = 0;
  ram[1219]  = 137;
  ram[1220]  = 255;
  ram[1221]  = 255;
  ram[1222]  = 255;
  ram[1223]  = 255;
  ram[1224]  = 255;
  ram[1225]  = 255;
  ram[1226]  = 255;
  ram[1227]  = 255;
  ram[1228]  = 255;
  ram[1229]  = 255;
  ram[1230]  = 255;
  ram[1231]  = 255;
  ram[1232]  = 255;
  ram[1233]  = 255;
  ram[1234]  = 255;
  ram[1235]  = 255;
  ram[1236]  = 255;
  ram[1237]  = 255;
  ram[1238]  = 71;
  ram[1239]  = 0;
  ram[1240]  = 0;
  ram[1241]  = 0;
  ram[1242]  = 0;
  ram[1243]  = 0;
  ram[1244]  = 0;
  ram[1245]  = 0;
  ram[1246]  = 0;
  ram[1247]  = 0;
  ram[1248]  = 0;
  ram[1249]  = 0;
  ram[1250]  = 0;
  ram[1251]  = 0;
  ram[1252]  = 0;
  ram[1253]  = 0;
  ram[1254]  = 0;
  ram[1255]  = 0;
  ram[1256]  = 0;
  ram[1257]  = 0;
  ram[1258]  = 0;
  ram[1259]  = 0;
  ram[1260]  = 0;
  ram[1261]  = 71;
  ram[1262]  = 255;
  ram[1263]  = 255;
  ram[1264]  = 255;
  ram[1265]  = 255;
  ram[1266]  = 255;
  ram[1267]  = 255;
  ram[1268]  = 255;
  ram[1269]  = 255;
  ram[1270]  = 255;
  ram[1271]  = 255;
  ram[1272]  = 255;
  ram[1273]  = 255;
  ram[1274]  = 255;
  ram[1275]  = 71;
  ram[1276]  = 0;
  ram[1277]  = 195;
  ram[1278]  = 255;
  ram[1279]  = 255;
  ram[1280]  = 255;
  ram[1281]  = 255;
  ram[1282]  = 255;
  ram[1283]  = 255;
  ram[1284]  = 255;
  ram[1285]  = 255;
  ram[1286]  = 105;
  ram[1287]  = 0;
  ram[1288]  = 71;
  ram[1289]  = 255;
  ram[1290]  = 255;
  ram[1291]  = 255;
  ram[1292]  = 255;
  ram[1293]  = 255;
  ram[1294]  = 255;
  ram[1295]  = 255;
  ram[1296]  = 255;
  ram[1297]  = 255;
  ram[1298]  = 255;
  ram[1299]  = 255;
  ram[1300]  = 255;
  ram[1301]  = 255;
  ram[1302]  = 255;
  ram[1303]  = 255;
  ram[1304]  = 255;
  ram[1305]  = 255;
  ram[1306]  = 255;
  ram[1307]  = 255;
  ram[1308]  = 255;
  ram[1309]  = 255;
  ram[1310]  = 255;
  ram[1311]  = 255;
  ram[1312]  = 255;
  ram[1313]  = 255;
  ram[1314]  = 255;
  ram[1315]  = 255;
  ram[1316]  = 255;
  ram[1317]  = 255;
  ram[1318]  = 255;
  ram[1319]  = 255;
  ram[1320]  = 255;
  ram[1321]  = 255;
  ram[1322]  = 255;
  ram[1323]  = 255;
  ram[1324]  = 255;
  ram[1325]  = 255;
  ram[1326]  = 255;
  ram[1327]  = 236;
  ram[1328]  = 52;
  ram[1329]  = 0;
  ram[1330]  = 0;
  ram[1331]  = 0;
  ram[1332]  = 35;
  ram[1333]  = 71;
  ram[1334]  = 122;
  ram[1335]  = 105;
  ram[1336]  = 71;
  ram[1337]  = 17;
  ram[1338]  = 0;
  ram[1339]  = 137;
  ram[1340]  = 255;
  ram[1341]  = 255;
  ram[1342]  = 255;
  ram[1343]  = 255;
  ram[1344]  = 255;
  ram[1345]  = 255;
  ram[1346]  = 255;
  ram[1347]  = 255;
  ram[1348]  = 255;
  ram[1349]  = 255;
  ram[1350]  = 255;
  ram[1351]  = 255;
  ram[1352]  = 255;
  ram[1353]  = 255;
  ram[1354]  = 255;
  ram[1355]  = 255;
  ram[1356]  = 255;
  ram[1357]  = 255;
  ram[1358]  = 167;
  ram[1359]  = 137;
  ram[1360]  = 137;
  ram[1361]  = 137;
  ram[1362]  = 137;
  ram[1363]  = 137;
  ram[1364]  = 0;
  ram[1365]  = 0;
  ram[1366]  = 137;
  ram[1367]  = 137;
  ram[1368]  = 137;
  ram[1369]  = 137;
  ram[1370]  = 137;
  ram[1371]  = 137;
  ram[1372]  = 137;
  ram[1373]  = 137;
  ram[1374]  = 35;
  ram[1375]  = 0;
  ram[1376]  = 71;
  ram[1377]  = 137;
  ram[1378]  = 137;
  ram[1379]  = 137;
  ram[1380]  = 137;
  ram[1381]  = 167;
  ram[1382]  = 255;
  ram[1383]  = 255;
  ram[1384]  = 255;
  ram[1385]  = 255;
  ram[1386]  = 255;
  ram[1387]  = 255;
  ram[1388]  = 255;
  ram[1389]  = 255;
  ram[1390]  = 255;
  ram[1391]  = 255;
  ram[1392]  = 255;
  ram[1393]  = 255;
  ram[1394]  = 255;
  ram[1395]  = 0;
  ram[1396]  = 0;
  ram[1397]  = 208;
  ram[1398]  = 255;
  ram[1399]  = 255;
  ram[1400]  = 255;
  ram[1401]  = 255;
  ram[1402]  = 255;
  ram[1403]  = 255;
  ram[1404]  = 255;
  ram[1405]  = 221;
  ram[1406]  = 0;
  ram[1407]  = 0;
  ram[1408]  = 195;
  ram[1409]  = 255;
  ram[1410]  = 255;
  ram[1411]  = 236;
  ram[1412]  = 137;
  ram[1413]  = 137;
  ram[1414]  = 255;
  ram[1415]  = 255;
  ram[1416]  = 255;
  ram[1417]  = 255;
  ram[1418]  = 255;
  ram[1419]  = 255;
  ram[1420]  = 255;
  ram[1421]  = 255;
  ram[1422]  = 255;
  ram[1423]  = 255;
  ram[1424]  = 255;
  ram[1425]  = 255;
  ram[1426]  = 255;
  ram[1427]  = 255;
  ram[1428]  = 255;
  ram[1429]  = 255;
  ram[1430]  = 255;
  ram[1431]  = 255;
  ram[1432]  = 255;
  ram[1433]  = 255;
  ram[1434]  = 255;
  ram[1435]  = 255;
  ram[1436]  = 255;
  ram[1437]  = 255;
  ram[1438]  = 255;
  ram[1439]  = 255;
  ram[1440]  = 255;
  ram[1441]  = 255;
  ram[1442]  = 255;
  ram[1443]  = 255;
  ram[1444]  = 255;
  ram[1445]  = 255;
  ram[1446]  = 236;
  ram[1447]  = 52;
  ram[1448]  = 0;
  ram[1449]  = 0;
  ram[1450]  = 52;
  ram[1451]  = 195;
  ram[1452]  = 255;
  ram[1453]  = 255;
  ram[1454]  = 255;
  ram[1455]  = 255;
  ram[1456]  = 255;
  ram[1457]  = 255;
  ram[1458]  = 181;
  ram[1459]  = 181;
  ram[1460]  = 255;
  ram[1461]  = 255;
  ram[1462]  = 255;
  ram[1463]  = 255;
  ram[1464]  = 255;
  ram[1465]  = 255;
  ram[1466]  = 255;
  ram[1467]  = 255;
  ram[1468]  = 255;
  ram[1469]  = 255;
  ram[1470]  = 255;
  ram[1471]  = 255;
  ram[1472]  = 255;
  ram[1473]  = 255;
  ram[1474]  = 255;
  ram[1475]  = 255;
  ram[1476]  = 255;
  ram[1477]  = 255;
  ram[1478]  = 255;
  ram[1479]  = 255;
  ram[1480]  = 255;
  ram[1481]  = 255;
  ram[1482]  = 255;
  ram[1483]  = 255;
  ram[1484]  = 0;
  ram[1485]  = 0;
  ram[1486]  = 255;
  ram[1487]  = 255;
  ram[1488]  = 255;
  ram[1489]  = 255;
  ram[1490]  = 255;
  ram[1491]  = 255;
  ram[1492]  = 255;
  ram[1493]  = 255;
  ram[1494]  = 71;
  ram[1495]  = 0;
  ram[1496]  = 137;
  ram[1497]  = 255;
  ram[1498]  = 255;
  ram[1499]  = 255;
  ram[1500]  = 255;
  ram[1501]  = 255;
  ram[1502]  = 255;
  ram[1503]  = 255;
  ram[1504]  = 255;
  ram[1505]  = 255;
  ram[1506]  = 255;
  ram[1507]  = 255;
  ram[1508]  = 255;
  ram[1509]  = 255;
  ram[1510]  = 255;
  ram[1511]  = 255;
  ram[1512]  = 255;
  ram[1513]  = 255;
  ram[1514]  = 221;
  ram[1515]  = 0;
  ram[1516]  = 0;
  ram[1517]  = 255;
  ram[1518]  = 255;
  ram[1519]  = 255;
  ram[1520]  = 255;
  ram[1521]  = 255;
  ram[1522]  = 255;
  ram[1523]  = 255;
  ram[1524]  = 255;
  ram[1525]  = 105;
  ram[1526]  = 0;
  ram[1527]  = 87;
  ram[1528]  = 255;
  ram[1529]  = 255;
  ram[1530]  = 255;
  ram[1531]  = 221;
  ram[1532]  = 0;
  ram[1533]  = 0;
  ram[1534]  = 208;
  ram[1535]  = 255;
  ram[1536]  = 255;
  ram[1537]  = 255;
  ram[1538]  = 255;
  ram[1539]  = 255;
  ram[1540]  = 255;
  ram[1541]  = 255;
  ram[1542]  = 255;
  ram[1543]  = 255;
  ram[1544]  = 255;
  ram[1545]  = 255;
  ram[1546]  = 255;
  ram[1547]  = 255;
  ram[1548]  = 255;
  ram[1549]  = 255;
  ram[1550]  = 255;
  ram[1551]  = 255;
  ram[1552]  = 255;
  ram[1553]  = 255;
  ram[1554]  = 255;
  ram[1555]  = 255;
  ram[1556]  = 255;
  ram[1557]  = 255;
  ram[1558]  = 255;
  ram[1559]  = 255;
  ram[1560]  = 255;
  ram[1561]  = 255;
  ram[1562]  = 255;
  ram[1563]  = 255;
  ram[1564]  = 255;
  ram[1565]  = 255;
  ram[1566]  = 71;
  ram[1567]  = 0;
  ram[1568]  = 0;
  ram[1569]  = 105;
  ram[1570]  = 255;
  ram[1571]  = 255;
  ram[1572]  = 255;
  ram[1573]  = 255;
  ram[1574]  = 255;
  ram[1575]  = 255;
  ram[1576]  = 255;
  ram[1577]  = 255;
  ram[1578]  = 255;
  ram[1579]  = 255;
  ram[1580]  = 255;
  ram[1581]  = 255;
  ram[1582]  = 255;
  ram[1583]  = 255;
  ram[1584]  = 255;
  ram[1585]  = 255;
  ram[1586]  = 255;
  ram[1587]  = 255;
  ram[1588]  = 255;
  ram[1589]  = 255;
  ram[1590]  = 255;
  ram[1591]  = 255;
  ram[1592]  = 255;
  ram[1593]  = 255;
  ram[1594]  = 255;
  ram[1595]  = 255;
  ram[1596]  = 255;
  ram[1597]  = 255;
  ram[1598]  = 255;
  ram[1599]  = 255;
  ram[1600]  = 255;
  ram[1601]  = 255;
  ram[1602]  = 255;
  ram[1603]  = 255;
  ram[1604]  = 0;
  ram[1605]  = 0;
  ram[1606]  = 255;
  ram[1607]  = 255;
  ram[1608]  = 255;
  ram[1609]  = 255;
  ram[1610]  = 255;
  ram[1611]  = 255;
  ram[1612]  = 255;
  ram[1613]  = 255;
  ram[1614]  = 71;
  ram[1615]  = 0;
  ram[1616]  = 137;
  ram[1617]  = 255;
  ram[1618]  = 255;
  ram[1619]  = 255;
  ram[1620]  = 255;
  ram[1621]  = 255;
  ram[1622]  = 255;
  ram[1623]  = 255;
  ram[1624]  = 255;
  ram[1625]  = 255;
  ram[1626]  = 255;
  ram[1627]  = 255;
  ram[1628]  = 255;
  ram[1629]  = 255;
  ram[1630]  = 255;
  ram[1631]  = 208;
  ram[1632]  = 71;
  ram[1633]  = 71;
  ram[1634]  = 52;
  ram[1635]  = 0;
  ram[1636]  = 17;
  ram[1637]  = 71;
  ram[1638]  = 71;
  ram[1639]  = 71;
  ram[1640]  = 71;
  ram[1641]  = 122;
  ram[1642]  = 255;
  ram[1643]  = 255;
  ram[1644]  = 208;
  ram[1645]  = 0;
  ram[1646]  = 0;
  ram[1647]  = 221;
  ram[1648]  = 255;
  ram[1649]  = 255;
  ram[1650]  = 255;
  ram[1651]  = 255;
  ram[1652]  = 137;
  ram[1653]  = 0;
  ram[1654]  = 71;
  ram[1655]  = 255;
  ram[1656]  = 255;
  ram[1657]  = 255;
  ram[1658]  = 255;
  ram[1659]  = 255;
  ram[1660]  = 255;
  ram[1661]  = 255;
  ram[1662]  = 255;
  ram[1663]  = 255;
  ram[1664]  = 255;
  ram[1665]  = 255;
  ram[1666]  = 255;
  ram[1667]  = 255;
  ram[1668]  = 255;
  ram[1669]  = 255;
  ram[1670]  = 255;
  ram[1671]  = 255;
  ram[1672]  = 255;
  ram[1673]  = 255;
  ram[1674]  = 255;
  ram[1675]  = 255;
  ram[1676]  = 255;
  ram[1677]  = 255;
  ram[1678]  = 255;
  ram[1679]  = 255;
  ram[1680]  = 255;
  ram[1681]  = 255;
  ram[1682]  = 255;
  ram[1683]  = 255;
  ram[1684]  = 255;
  ram[1685]  = 167;
  ram[1686]  = 0;
  ram[1687]  = 0;
  ram[1688]  = 71;
  ram[1689]  = 255;
  ram[1690]  = 255;
  ram[1691]  = 255;
  ram[1692]  = 255;
  ram[1693]  = 255;
  ram[1694]  = 255;
  ram[1695]  = 255;
  ram[1696]  = 255;
  ram[1697]  = 255;
  ram[1698]  = 255;
  ram[1699]  = 255;
  ram[1700]  = 255;
  ram[1701]  = 255;
  ram[1702]  = 255;
  ram[1703]  = 255;
  ram[1704]  = 255;
  ram[1705]  = 255;
  ram[1706]  = 255;
  ram[1707]  = 255;
  ram[1708]  = 255;
  ram[1709]  = 255;
  ram[1710]  = 255;
  ram[1711]  = 255;
  ram[1712]  = 255;
  ram[1713]  = 255;
  ram[1714]  = 255;
  ram[1715]  = 255;
  ram[1716]  = 255;
  ram[1717]  = 255;
  ram[1718]  = 255;
  ram[1719]  = 255;
  ram[1720]  = 255;
  ram[1721]  = 255;
  ram[1722]  = 255;
  ram[1723]  = 255;
  ram[1724]  = 0;
  ram[1725]  = 0;
  ram[1726]  = 255;
  ram[1727]  = 255;
  ram[1728]  = 255;
  ram[1729]  = 255;
  ram[1730]  = 255;
  ram[1731]  = 255;
  ram[1732]  = 255;
  ram[1733]  = 255;
  ram[1734]  = 71;
  ram[1735]  = 0;
  ram[1736]  = 137;
  ram[1737]  = 255;
  ram[1738]  = 255;
  ram[1739]  = 255;
  ram[1740]  = 255;
  ram[1741]  = 255;
  ram[1742]  = 255;
  ram[1743]  = 255;
  ram[1744]  = 255;
  ram[1745]  = 255;
  ram[1746]  = 255;
  ram[1747]  = 255;
  ram[1748]  = 255;
  ram[1749]  = 255;
  ram[1750]  = 255;
  ram[1751]  = 195;
  ram[1752]  = 0;
  ram[1753]  = 0;
  ram[1754]  = 0;
  ram[1755]  = 0;
  ram[1756]  = 0;
  ram[1757]  = 0;
  ram[1758]  = 0;
  ram[1759]  = 0;
  ram[1760]  = 0;
  ram[1761]  = 71;
  ram[1762]  = 255;
  ram[1763]  = 255;
  ram[1764]  = 71;
  ram[1765]  = 0;
  ram[1766]  = 137;
  ram[1767]  = 255;
  ram[1768]  = 255;
  ram[1769]  = 255;
  ram[1770]  = 255;
  ram[1771]  = 255;
  ram[1772]  = 236;
  ram[1773]  = 17;
  ram[1774]  = 0;
  ram[1775]  = 167;
  ram[1776]  = 255;
  ram[1777]  = 255;
  ram[1778]  = 255;
  ram[1779]  = 255;
  ram[1780]  = 255;
  ram[1781]  = 255;
  ram[1782]  = 255;
  ram[1783]  = 255;
  ram[1784]  = 255;
  ram[1785]  = 255;
  ram[1786]  = 255;
  ram[1787]  = 255;
  ram[1788]  = 255;
  ram[1789]  = 255;
  ram[1790]  = 255;
  ram[1791]  = 255;
  ram[1792]  = 255;
  ram[1793]  = 255;
  ram[1794]  = 255;
  ram[1795]  = 255;
  ram[1796]  = 255;
  ram[1797]  = 255;
  ram[1798]  = 255;
  ram[1799]  = 255;
  ram[1800]  = 255;
  ram[1801]  = 255;
  ram[1802]  = 255;
  ram[1803]  = 255;
  ram[1804]  = 255;
  ram[1805]  = 35;
  ram[1806]  = 0;
  ram[1807]  = 0;
  ram[1808]  = 221;
  ram[1809]  = 255;
  ram[1810]  = 255;
  ram[1811]  = 255;
  ram[1812]  = 255;
  ram[1813]  = 255;
  ram[1814]  = 255;
  ram[1815]  = 255;
  ram[1816]  = 255;
  ram[1817]  = 255;
  ram[1818]  = 255;
  ram[1819]  = 255;
  ram[1820]  = 255;
  ram[1821]  = 255;
  ram[1822]  = 255;
  ram[1823]  = 255;
  ram[1824]  = 255;
  ram[1825]  = 255;
  ram[1826]  = 255;
  ram[1827]  = 255;
  ram[1828]  = 255;
  ram[1829]  = 255;
  ram[1830]  = 255;
  ram[1831]  = 255;
  ram[1832]  = 255;
  ram[1833]  = 255;
  ram[1834]  = 255;
  ram[1835]  = 255;
  ram[1836]  = 255;
  ram[1837]  = 255;
  ram[1838]  = 255;
  ram[1839]  = 255;
  ram[1840]  = 255;
  ram[1841]  = 255;
  ram[1842]  = 255;
  ram[1843]  = 255;
  ram[1844]  = 0;
  ram[1845]  = 0;
  ram[1846]  = 255;
  ram[1847]  = 255;
  ram[1848]  = 255;
  ram[1849]  = 255;
  ram[1850]  = 255;
  ram[1851]  = 255;
  ram[1852]  = 255;
  ram[1853]  = 255;
  ram[1854]  = 71;
  ram[1855]  = 0;
  ram[1856]  = 137;
  ram[1857]  = 255;
  ram[1858]  = 255;
  ram[1859]  = 255;
  ram[1860]  = 255;
  ram[1861]  = 255;
  ram[1862]  = 255;
  ram[1863]  = 255;
  ram[1864]  = 255;
  ram[1865]  = 255;
  ram[1866]  = 255;
  ram[1867]  = 255;
  ram[1868]  = 255;
  ram[1869]  = 255;
  ram[1870]  = 255;
  ram[1871]  = 236;
  ram[1872]  = 195;
  ram[1873]  = 195;
  ram[1874]  = 71;
  ram[1875]  = 0;
  ram[1876]  = 122;
  ram[1877]  = 195;
  ram[1878]  = 195;
  ram[1879]  = 152;
  ram[1880]  = 0;
  ram[1881]  = 71;
  ram[1882]  = 255;
  ram[1883]  = 152;
  ram[1884]  = 0;
  ram[1885]  = 35;
  ram[1886]  = 236;
  ram[1887]  = 255;
  ram[1888]  = 255;
  ram[1889]  = 255;
  ram[1890]  = 255;
  ram[1891]  = 255;
  ram[1892]  = 255;
  ram[1893]  = 137;
  ram[1894]  = 0;
  ram[1895]  = 35;
  ram[1896]  = 236;
  ram[1897]  = 255;
  ram[1898]  = 255;
  ram[1899]  = 255;
  ram[1900]  = 255;
  ram[1901]  = 255;
  ram[1902]  = 255;
  ram[1903]  = 255;
  ram[1904]  = 255;
  ram[1905]  = 255;
  ram[1906]  = 255;
  ram[1907]  = 255;
  ram[1908]  = 255;
  ram[1909]  = 255;
  ram[1910]  = 255;
  ram[1911]  = 255;
  ram[1912]  = 255;
  ram[1913]  = 255;
  ram[1914]  = 255;
  ram[1915]  = 255;
  ram[1916]  = 255;
  ram[1917]  = 255;
  ram[1918]  = 255;
  ram[1919]  = 255;
  ram[1920]  = 255;
  ram[1921]  = 255;
  ram[1922]  = 255;
  ram[1923]  = 255;
  ram[1924]  = 208;
  ram[1925]  = 0;
  ram[1926]  = 0;
  ram[1927]  = 105;
  ram[1928]  = 255;
  ram[1929]  = 255;
  ram[1930]  = 255;
  ram[1931]  = 255;
  ram[1932]  = 255;
  ram[1933]  = 255;
  ram[1934]  = 255;
  ram[1935]  = 255;
  ram[1936]  = 255;
  ram[1937]  = 255;
  ram[1938]  = 255;
  ram[1939]  = 255;
  ram[1940]  = 255;
  ram[1941]  = 255;
  ram[1942]  = 255;
  ram[1943]  = 255;
  ram[1944]  = 255;
  ram[1945]  = 255;
  ram[1946]  = 255;
  ram[1947]  = 255;
  ram[1948]  = 255;
  ram[1949]  = 255;
  ram[1950]  = 255;
  ram[1951]  = 255;
  ram[1952]  = 255;
  ram[1953]  = 255;
  ram[1954]  = 255;
  ram[1955]  = 255;
  ram[1956]  = 255;
  ram[1957]  = 255;
  ram[1958]  = 255;
  ram[1959]  = 255;
  ram[1960]  = 255;
  ram[1961]  = 255;
  ram[1962]  = 255;
  ram[1963]  = 255;
  ram[1964]  = 0;
  ram[1965]  = 0;
  ram[1966]  = 255;
  ram[1967]  = 255;
  ram[1968]  = 255;
  ram[1969]  = 255;
  ram[1970]  = 255;
  ram[1971]  = 255;
  ram[1972]  = 255;
  ram[1973]  = 255;
  ram[1974]  = 71;
  ram[1975]  = 0;
  ram[1976]  = 137;
  ram[1977]  = 255;
  ram[1978]  = 255;
  ram[1979]  = 255;
  ram[1980]  = 255;
  ram[1981]  = 255;
  ram[1982]  = 255;
  ram[1983]  = 255;
  ram[1984]  = 255;
  ram[1985]  = 255;
  ram[1986]  = 255;
  ram[1987]  = 255;
  ram[1988]  = 255;
  ram[1989]  = 255;
  ram[1990]  = 255;
  ram[1991]  = 255;
  ram[1992]  = 255;
  ram[1993]  = 255;
  ram[1994]  = 71;
  ram[1995]  = 0;
  ram[1996]  = 195;
  ram[1997]  = 255;
  ram[1998]  = 255;
  ram[1999]  = 167;
  ram[2000]  = 0;
  ram[2001]  = 105;
  ram[2002]  = 195;
  ram[2003]  = 17;
  ram[2004]  = 0;
  ram[2005]  = 87;
  ram[2006]  = 137;
  ram[2007]  = 137;
  ram[2008]  = 71;
  ram[2009]  = 71;
  ram[2010]  = 71;
  ram[2011]  = 71;
  ram[2012]  = 17;
  ram[2013]  = 0;
  ram[2014]  = 0;
  ram[2015]  = 0;
  ram[2016]  = 137;
  ram[2017]  = 255;
  ram[2018]  = 255;
  ram[2019]  = 255;
  ram[2020]  = 255;
  ram[2021]  = 255;
  ram[2022]  = 255;
  ram[2023]  = 255;
  ram[2024]  = 255;
  ram[2025]  = 255;
  ram[2026]  = 255;
  ram[2027]  = 255;
  ram[2028]  = 255;
  ram[2029]  = 255;
  ram[2030]  = 255;
  ram[2031]  = 255;
  ram[2032]  = 255;
  ram[2033]  = 255;
  ram[2034]  = 255;
  ram[2035]  = 255;
  ram[2036]  = 255;
  ram[2037]  = 255;
  ram[2038]  = 255;
  ram[2039]  = 255;
  ram[2040]  = 255;
  ram[2041]  = 255;
  ram[2042]  = 255;
  ram[2043]  = 255;
  ram[2044]  = 152;
  ram[2045]  = 0;
  ram[2046]  = 0;
  ram[2047]  = 167;
  ram[2048]  = 255;
  ram[2049]  = 255;
  ram[2050]  = 255;
  ram[2051]  = 255;
  ram[2052]  = 255;
  ram[2053]  = 255;
  ram[2054]  = 255;
  ram[2055]  = 255;
  ram[2056]  = 255;
  ram[2057]  = 255;
  ram[2058]  = 255;
  ram[2059]  = 255;
  ram[2060]  = 255;
  ram[2061]  = 255;
  ram[2062]  = 255;
  ram[2063]  = 255;
  ram[2064]  = 255;
  ram[2065]  = 255;
  ram[2066]  = 255;
  ram[2067]  = 255;
  ram[2068]  = 255;
  ram[2069]  = 255;
  ram[2070]  = 255;
  ram[2071]  = 255;
  ram[2072]  = 255;
  ram[2073]  = 255;
  ram[2074]  = 255;
  ram[2075]  = 255;
  ram[2076]  = 255;
  ram[2077]  = 255;
  ram[2078]  = 255;
  ram[2079]  = 255;
  ram[2080]  = 255;
  ram[2081]  = 255;
  ram[2082]  = 255;
  ram[2083]  = 255;
  ram[2084]  = 0;
  ram[2085]  = 0;
  ram[2086]  = 255;
  ram[2087]  = 255;
  ram[2088]  = 255;
  ram[2089]  = 255;
  ram[2090]  = 255;
  ram[2091]  = 255;
  ram[2092]  = 255;
  ram[2093]  = 255;
  ram[2094]  = 71;
  ram[2095]  = 0;
  ram[2096]  = 137;
  ram[2097]  = 255;
  ram[2098]  = 255;
  ram[2099]  = 255;
  ram[2100]  = 255;
  ram[2101]  = 255;
  ram[2102]  = 255;
  ram[2103]  = 255;
  ram[2104]  = 255;
  ram[2105]  = 255;
  ram[2106]  = 255;
  ram[2107]  = 255;
  ram[2108]  = 255;
  ram[2109]  = 255;
  ram[2110]  = 255;
  ram[2111]  = 255;
  ram[2112]  = 255;
  ram[2113]  = 255;
  ram[2114]  = 0;
  ram[2115]  = 0;
  ram[2116]  = 255;
  ram[2117]  = 255;
  ram[2118]  = 255;
  ram[2119]  = 137;
  ram[2120]  = 0;
  ram[2121]  = 137;
  ram[2122]  = 35;
  ram[2123]  = 0;
  ram[2124]  = 0;
  ram[2125]  = 0;
  ram[2126]  = 0;
  ram[2127]  = 0;
  ram[2128]  = 0;
  ram[2129]  = 0;
  ram[2130]  = 0;
  ram[2131]  = 0;
  ram[2132]  = 0;
  ram[2133]  = 0;
  ram[2134]  = 52;
  ram[2135]  = 0;
  ram[2136]  = 17;
  ram[2137]  = 236;
  ram[2138]  = 255;
  ram[2139]  = 255;
  ram[2140]  = 255;
  ram[2141]  = 255;
  ram[2142]  = 255;
  ram[2143]  = 255;
  ram[2144]  = 255;
  ram[2145]  = 255;
  ram[2146]  = 255;
  ram[2147]  = 255;
  ram[2148]  = 255;
  ram[2149]  = 255;
  ram[2150]  = 255;
  ram[2151]  = 255;
  ram[2152]  = 255;
  ram[2153]  = 255;
  ram[2154]  = 255;
  ram[2155]  = 255;
  ram[2156]  = 255;
  ram[2157]  = 255;
  ram[2158]  = 255;
  ram[2159]  = 255;
  ram[2160]  = 255;
  ram[2161]  = 255;
  ram[2162]  = 255;
  ram[2163]  = 255;
  ram[2164]  = 122;
  ram[2165]  = 0;
  ram[2166]  = 0;
  ram[2167]  = 195;
  ram[2168]  = 255;
  ram[2169]  = 255;
  ram[2170]  = 255;
  ram[2171]  = 255;
  ram[2172]  = 255;
  ram[2173]  = 255;
  ram[2174]  = 255;
  ram[2175]  = 255;
  ram[2176]  = 255;
  ram[2177]  = 255;
  ram[2178]  = 255;
  ram[2179]  = 255;
  ram[2180]  = 255;
  ram[2181]  = 255;
  ram[2182]  = 255;
  ram[2183]  = 255;
  ram[2184]  = 255;
  ram[2185]  = 255;
  ram[2186]  = 255;
  ram[2187]  = 255;
  ram[2188]  = 255;
  ram[2189]  = 255;
  ram[2190]  = 255;
  ram[2191]  = 255;
  ram[2192]  = 255;
  ram[2193]  = 255;
  ram[2194]  = 255;
  ram[2195]  = 255;
  ram[2196]  = 255;
  ram[2197]  = 255;
  ram[2198]  = 255;
  ram[2199]  = 255;
  ram[2200]  = 255;
  ram[2201]  = 255;
  ram[2202]  = 255;
  ram[2203]  = 255;
  ram[2204]  = 0;
  ram[2205]  = 0;
  ram[2206]  = 255;
  ram[2207]  = 255;
  ram[2208]  = 255;
  ram[2209]  = 255;
  ram[2210]  = 255;
  ram[2211]  = 255;
  ram[2212]  = 255;
  ram[2213]  = 255;
  ram[2214]  = 71;
  ram[2215]  = 0;
  ram[2216]  = 137;
  ram[2217]  = 255;
  ram[2218]  = 255;
  ram[2219]  = 255;
  ram[2220]  = 255;
  ram[2221]  = 255;
  ram[2222]  = 255;
  ram[2223]  = 255;
  ram[2224]  = 255;
  ram[2225]  = 255;
  ram[2226]  = 255;
  ram[2227]  = 255;
  ram[2228]  = 255;
  ram[2229]  = 255;
  ram[2230]  = 255;
  ram[2231]  = 255;
  ram[2232]  = 255;
  ram[2233]  = 208;
  ram[2234]  = 0;
  ram[2235]  = 52;
  ram[2236]  = 255;
  ram[2237]  = 255;
  ram[2238]  = 255;
  ram[2239]  = 105;
  ram[2240]  = 0;
  ram[2241]  = 167;
  ram[2242]  = 167;
  ram[2243]  = 35;
  ram[2244]  = 87;
  ram[2245]  = 137;
  ram[2246]  = 137;
  ram[2247]  = 167;
  ram[2248]  = 195;
  ram[2249]  = 195;
  ram[2250]  = 221;
  ram[2251]  = 255;
  ram[2252]  = 255;
  ram[2253]  = 255;
  ram[2254]  = 236;
  ram[2255]  = 17;
  ram[2256]  = 0;
  ram[2257]  = 137;
  ram[2258]  = 255;
  ram[2259]  = 255;
  ram[2260]  = 255;
  ram[2261]  = 255;
  ram[2262]  = 255;
  ram[2263]  = 255;
  ram[2264]  = 255;
  ram[2265]  = 255;
  ram[2266]  = 255;
  ram[2267]  = 255;
  ram[2268]  = 255;
  ram[2269]  = 255;
  ram[2270]  = 255;
  ram[2271]  = 255;
  ram[2272]  = 255;
  ram[2273]  = 255;
  ram[2274]  = 255;
  ram[2275]  = 255;
  ram[2276]  = 255;
  ram[2277]  = 255;
  ram[2278]  = 255;
  ram[2279]  = 255;
  ram[2280]  = 255;
  ram[2281]  = 255;
  ram[2282]  = 255;
  ram[2283]  = 255;
  ram[2284]  = 71;
  ram[2285]  = 0;
  ram[2286]  = 0;
  ram[2287]  = 255;
  ram[2288]  = 255;
  ram[2289]  = 255;
  ram[2290]  = 255;
  ram[2291]  = 255;
  ram[2292]  = 255;
  ram[2293]  = 255;
  ram[2294]  = 255;
  ram[2295]  = 255;
  ram[2296]  = 255;
  ram[2297]  = 255;
  ram[2298]  = 255;
  ram[2299]  = 255;
  ram[2300]  = 255;
  ram[2301]  = 255;
  ram[2302]  = 255;
  ram[2303]  = 255;
  ram[2304]  = 255;
  ram[2305]  = 255;
  ram[2306]  = 255;
  ram[2307]  = 255;
  ram[2308]  = 255;
  ram[2309]  = 255;
  ram[2310]  = 255;
  ram[2311]  = 255;
  ram[2312]  = 255;
  ram[2313]  = 255;
  ram[2314]  = 255;
  ram[2315]  = 255;
  ram[2316]  = 255;
  ram[2317]  = 71;
  ram[2318]  = 71;
  ram[2319]  = 71;
  ram[2320]  = 71;
  ram[2321]  = 71;
  ram[2322]  = 71;
  ram[2323]  = 71;
  ram[2324]  = 0;
  ram[2325]  = 0;
  ram[2326]  = 71;
  ram[2327]  = 71;
  ram[2328]  = 71;
  ram[2329]  = 71;
  ram[2330]  = 71;
  ram[2331]  = 71;
  ram[2332]  = 71;
  ram[2333]  = 71;
  ram[2334]  = 17;
  ram[2335]  = 0;
  ram[2336]  = 35;
  ram[2337]  = 71;
  ram[2338]  = 71;
  ram[2339]  = 71;
  ram[2340]  = 71;
  ram[2341]  = 71;
  ram[2342]  = 71;
  ram[2343]  = 255;
  ram[2344]  = 255;
  ram[2345]  = 255;
  ram[2346]  = 255;
  ram[2347]  = 255;
  ram[2348]  = 255;
  ram[2349]  = 255;
  ram[2350]  = 255;
  ram[2351]  = 255;
  ram[2352]  = 255;
  ram[2353]  = 167;
  ram[2354]  = 0;
  ram[2355]  = 105;
  ram[2356]  = 255;
  ram[2357]  = 255;
  ram[2358]  = 255;
  ram[2359]  = 71;
  ram[2360]  = 0;
  ram[2361]  = 208;
  ram[2362]  = 255;
  ram[2363]  = 255;
  ram[2364]  = 255;
  ram[2365]  = 255;
  ram[2366]  = 255;
  ram[2367]  = 255;
  ram[2368]  = 255;
  ram[2369]  = 255;
  ram[2370]  = 255;
  ram[2371]  = 255;
  ram[2372]  = 255;
  ram[2373]  = 255;
  ram[2374]  = 255;
  ram[2375]  = 137;
  ram[2376]  = 17;
  ram[2377]  = 137;
  ram[2378]  = 255;
  ram[2379]  = 255;
  ram[2380]  = 255;
  ram[2381]  = 255;
  ram[2382]  = 255;
  ram[2383]  = 255;
  ram[2384]  = 255;
  ram[2385]  = 255;
  ram[2386]  = 255;
  ram[2387]  = 255;
  ram[2388]  = 255;
  ram[2389]  = 255;
  ram[2390]  = 255;
  ram[2391]  = 255;
  ram[2392]  = 255;
  ram[2393]  = 255;
  ram[2394]  = 255;
  ram[2395]  = 255;
  ram[2396]  = 255;
  ram[2397]  = 255;
  ram[2398]  = 255;
  ram[2399]  = 255;
  ram[2400]  = 255;
  ram[2401]  = 255;
  ram[2402]  = 255;
  ram[2403]  = 255;
  ram[2404]  = 71;
  ram[2405]  = 0;
  ram[2406]  = 0;
  ram[2407]  = 255;
  ram[2408]  = 255;
  ram[2409]  = 255;
  ram[2410]  = 255;
  ram[2411]  = 255;
  ram[2412]  = 255;
  ram[2413]  = 255;
  ram[2414]  = 255;
  ram[2415]  = 255;
  ram[2416]  = 255;
  ram[2417]  = 255;
  ram[2418]  = 255;
  ram[2419]  = 255;
  ram[2420]  = 255;
  ram[2421]  = 255;
  ram[2422]  = 255;
  ram[2423]  = 255;
  ram[2424]  = 255;
  ram[2425]  = 255;
  ram[2426]  = 255;
  ram[2427]  = 255;
  ram[2428]  = 255;
  ram[2429]  = 255;
  ram[2430]  = 255;
  ram[2431]  = 255;
  ram[2432]  = 255;
  ram[2433]  = 255;
  ram[2434]  = 255;
  ram[2435]  = 255;
  ram[2436]  = 255;
  ram[2437]  = 0;
  ram[2438]  = 0;
  ram[2439]  = 0;
  ram[2440]  = 0;
  ram[2441]  = 0;
  ram[2442]  = 0;
  ram[2443]  = 0;
  ram[2444]  = 0;
  ram[2445]  = 0;
  ram[2446]  = 0;
  ram[2447]  = 0;
  ram[2448]  = 0;
  ram[2449]  = 0;
  ram[2450]  = 0;
  ram[2451]  = 0;
  ram[2452]  = 0;
  ram[2453]  = 0;
  ram[2454]  = 0;
  ram[2455]  = 0;
  ram[2456]  = 0;
  ram[2457]  = 0;
  ram[2458]  = 0;
  ram[2459]  = 0;
  ram[2460]  = 0;
  ram[2461]  = 0;
  ram[2462]  = 0;
  ram[2463]  = 255;
  ram[2464]  = 255;
  ram[2465]  = 255;
  ram[2466]  = 255;
  ram[2467]  = 255;
  ram[2468]  = 255;
  ram[2469]  = 255;
  ram[2470]  = 255;
  ram[2471]  = 255;
  ram[2472]  = 255;
  ram[2473]  = 105;
  ram[2474]  = 0;
  ram[2475]  = 167;
  ram[2476]  = 255;
  ram[2477]  = 255;
  ram[2478]  = 255;
  ram[2479]  = 0;
  ram[2480]  = 0;
  ram[2481]  = 255;
  ram[2482]  = 255;
  ram[2483]  = 255;
  ram[2484]  = 255;
  ram[2485]  = 255;
  ram[2486]  = 255;
  ram[2487]  = 255;
  ram[2488]  = 255;
  ram[2489]  = 255;
  ram[2490]  = 255;
  ram[2491]  = 255;
  ram[2492]  = 255;
  ram[2493]  = 255;
  ram[2494]  = 255;
  ram[2495]  = 236;
  ram[2496]  = 236;
  ram[2497]  = 255;
  ram[2498]  = 255;
  ram[2499]  = 255;
  ram[2500]  = 255;
  ram[2501]  = 255;
  ram[2502]  = 255;
  ram[2503]  = 255;
  ram[2504]  = 255;
  ram[2505]  = 255;
  ram[2506]  = 255;
  ram[2507]  = 255;
  ram[2508]  = 255;
  ram[2509]  = 255;
  ram[2510]  = 255;
  ram[2511]  = 255;
  ram[2512]  = 255;
  ram[2513]  = 255;
  ram[2514]  = 255;
  ram[2515]  = 255;
  ram[2516]  = 255;
  ram[2517]  = 255;
  ram[2518]  = 255;
  ram[2519]  = 255;
  ram[2520]  = 255;
  ram[2521]  = 255;
  ram[2522]  = 255;
  ram[2523]  = 255;
  ram[2524]  = 105;
  ram[2525]  = 0;
  ram[2526]  = 0;
  ram[2527]  = 195;
  ram[2528]  = 255;
  ram[2529]  = 255;
  ram[2530]  = 255;
  ram[2531]  = 255;
  ram[2532]  = 255;
  ram[2533]  = 255;
  ram[2534]  = 255;
  ram[2535]  = 255;
  ram[2536]  = 255;
  ram[2537]  = 255;
  ram[2538]  = 255;
  ram[2539]  = 255;
  ram[2540]  = 255;
  ram[2541]  = 255;
  ram[2542]  = 255;
  ram[2543]  = 255;
  ram[2544]  = 255;
  ram[2545]  = 255;
  ram[2546]  = 255;
  ram[2547]  = 255;
  ram[2548]  = 255;
  ram[2549]  = 255;
  ram[2550]  = 255;
  ram[2551]  = 255;
  ram[2552]  = 255;
  ram[2553]  = 255;
  ram[2554]  = 255;
  ram[2555]  = 255;
  ram[2556]  = 255;
  ram[2557]  = 195;
  ram[2558]  = 195;
  ram[2559]  = 195;
  ram[2560]  = 195;
  ram[2561]  = 195;
  ram[2562]  = 195;
  ram[2563]  = 195;
  ram[2564]  = 0;
  ram[2565]  = 0;
  ram[2566]  = 195;
  ram[2567]  = 195;
  ram[2568]  = 195;
  ram[2569]  = 195;
  ram[2570]  = 195;
  ram[2571]  = 195;
  ram[2572]  = 195;
  ram[2573]  = 195;
  ram[2574]  = 52;
  ram[2575]  = 0;
  ram[2576]  = 105;
  ram[2577]  = 195;
  ram[2578]  = 195;
  ram[2579]  = 195;
  ram[2580]  = 195;
  ram[2581]  = 195;
  ram[2582]  = 195;
  ram[2583]  = 255;
  ram[2584]  = 255;
  ram[2585]  = 255;
  ram[2586]  = 255;
  ram[2587]  = 255;
  ram[2588]  = 255;
  ram[2589]  = 255;
  ram[2590]  = 255;
  ram[2591]  = 255;
  ram[2592]  = 255;
  ram[2593]  = 35;
  ram[2594]  = 0;
  ram[2595]  = 221;
  ram[2596]  = 255;
  ram[2597]  = 255;
  ram[2598]  = 195;
  ram[2599]  = 0;
  ram[2600]  = 71;
  ram[2601]  = 255;
  ram[2602]  = 255;
  ram[2603]  = 167;
  ram[2604]  = 137;
  ram[2605]  = 137;
  ram[2606]  = 137;
  ram[2607]  = 137;
  ram[2608]  = 137;
  ram[2609]  = 137;
  ram[2610]  = 137;
  ram[2611]  = 137;
  ram[2612]  = 137;
  ram[2613]  = 137;
  ram[2614]  = 137;
  ram[2615]  = 137;
  ram[2616]  = 255;
  ram[2617]  = 255;
  ram[2618]  = 255;
  ram[2619]  = 255;
  ram[2620]  = 255;
  ram[2621]  = 255;
  ram[2622]  = 255;
  ram[2623]  = 255;
  ram[2624]  = 255;
  ram[2625]  = 255;
  ram[2626]  = 255;
  ram[2627]  = 255;
  ram[2628]  = 255;
  ram[2629]  = 255;
  ram[2630]  = 255;
  ram[2631]  = 255;
  ram[2632]  = 255;
  ram[2633]  = 255;
  ram[2634]  = 255;
  ram[2635]  = 255;
  ram[2636]  = 255;
  ram[2637]  = 255;
  ram[2638]  = 255;
  ram[2639]  = 255;
  ram[2640]  = 255;
  ram[2641]  = 255;
  ram[2642]  = 255;
  ram[2643]  = 255;
  ram[2644]  = 137;
  ram[2645]  = 0;
  ram[2646]  = 0;
  ram[2647]  = 167;
  ram[2648]  = 255;
  ram[2649]  = 255;
  ram[2650]  = 255;
  ram[2651]  = 255;
  ram[2652]  = 255;
  ram[2653]  = 255;
  ram[2654]  = 255;
  ram[2655]  = 255;
  ram[2656]  = 255;
  ram[2657]  = 255;
  ram[2658]  = 255;
  ram[2659]  = 255;
  ram[2660]  = 255;
  ram[2661]  = 255;
  ram[2662]  = 255;
  ram[2663]  = 255;
  ram[2664]  = 255;
  ram[2665]  = 255;
  ram[2666]  = 255;
  ram[2667]  = 255;
  ram[2668]  = 255;
  ram[2669]  = 255;
  ram[2670]  = 255;
  ram[2671]  = 255;
  ram[2672]  = 255;
  ram[2673]  = 255;
  ram[2674]  = 255;
  ram[2675]  = 255;
  ram[2676]  = 255;
  ram[2677]  = 255;
  ram[2678]  = 255;
  ram[2679]  = 255;
  ram[2680]  = 255;
  ram[2681]  = 255;
  ram[2682]  = 255;
  ram[2683]  = 195;
  ram[2684]  = 0;
  ram[2685]  = 0;
  ram[2686]  = 255;
  ram[2687]  = 255;
  ram[2688]  = 255;
  ram[2689]  = 255;
  ram[2690]  = 255;
  ram[2691]  = 255;
  ram[2692]  = 255;
  ram[2693]  = 255;
  ram[2694]  = 71;
  ram[2695]  = 0;
  ram[2696]  = 137;
  ram[2697]  = 255;
  ram[2698]  = 255;
  ram[2699]  = 255;
  ram[2700]  = 255;
  ram[2701]  = 255;
  ram[2702]  = 255;
  ram[2703]  = 255;
  ram[2704]  = 255;
  ram[2705]  = 255;
  ram[2706]  = 255;
  ram[2707]  = 255;
  ram[2708]  = 255;
  ram[2709]  = 255;
  ram[2710]  = 255;
  ram[2711]  = 255;
  ram[2712]  = 236;
  ram[2713]  = 0;
  ram[2714]  = 0;
  ram[2715]  = 236;
  ram[2716]  = 255;
  ram[2717]  = 255;
  ram[2718]  = 122;
  ram[2719]  = 0;
  ram[2720]  = 137;
  ram[2721]  = 255;
  ram[2722]  = 255;
  ram[2723]  = 71;
  ram[2724]  = 0;
  ram[2725]  = 0;
  ram[2726]  = 0;
  ram[2727]  = 0;
  ram[2728]  = 0;
  ram[2729]  = 0;
  ram[2730]  = 0;
  ram[2731]  = 0;
  ram[2732]  = 0;
  ram[2733]  = 0;
  ram[2734]  = 0;
  ram[2735]  = 0;
  ram[2736]  = 255;
  ram[2737]  = 255;
  ram[2738]  = 255;
  ram[2739]  = 255;
  ram[2740]  = 255;
  ram[2741]  = 255;
  ram[2742]  = 255;
  ram[2743]  = 255;
  ram[2744]  = 255;
  ram[2745]  = 255;
  ram[2746]  = 255;
  ram[2747]  = 255;
  ram[2748]  = 255;
  ram[2749]  = 255;
  ram[2750]  = 255;
  ram[2751]  = 255;
  ram[2752]  = 255;
  ram[2753]  = 255;
  ram[2754]  = 255;
  ram[2755]  = 255;
  ram[2756]  = 255;
  ram[2757]  = 255;
  ram[2758]  = 255;
  ram[2759]  = 255;
  ram[2760]  = 255;
  ram[2761]  = 255;
  ram[2762]  = 255;
  ram[2763]  = 255;
  ram[2764]  = 181;
  ram[2765]  = 0;
  ram[2766]  = 0;
  ram[2767]  = 105;
  ram[2768]  = 255;
  ram[2769]  = 255;
  ram[2770]  = 255;
  ram[2771]  = 255;
  ram[2772]  = 255;
  ram[2773]  = 255;
  ram[2774]  = 255;
  ram[2775]  = 255;
  ram[2776]  = 255;
  ram[2777]  = 255;
  ram[2778]  = 255;
  ram[2779]  = 255;
  ram[2780]  = 255;
  ram[2781]  = 255;
  ram[2782]  = 255;
  ram[2783]  = 255;
  ram[2784]  = 255;
  ram[2785]  = 255;
  ram[2786]  = 255;
  ram[2787]  = 255;
  ram[2788]  = 255;
  ram[2789]  = 255;
  ram[2790]  = 255;
  ram[2791]  = 255;
  ram[2792]  = 255;
  ram[2793]  = 255;
  ram[2794]  = 255;
  ram[2795]  = 255;
  ram[2796]  = 255;
  ram[2797]  = 255;
  ram[2798]  = 255;
  ram[2799]  = 255;
  ram[2800]  = 255;
  ram[2801]  = 255;
  ram[2802]  = 255;
  ram[2803]  = 195;
  ram[2804]  = 0;
  ram[2805]  = 0;
  ram[2806]  = 255;
  ram[2807]  = 255;
  ram[2808]  = 255;
  ram[2809]  = 255;
  ram[2810]  = 255;
  ram[2811]  = 255;
  ram[2812]  = 255;
  ram[2813]  = 255;
  ram[2814]  = 71;
  ram[2815]  = 0;
  ram[2816]  = 137;
  ram[2817]  = 255;
  ram[2818]  = 255;
  ram[2819]  = 255;
  ram[2820]  = 255;
  ram[2821]  = 255;
  ram[2822]  = 255;
  ram[2823]  = 255;
  ram[2824]  = 255;
  ram[2825]  = 255;
  ram[2826]  = 255;
  ram[2827]  = 255;
  ram[2828]  = 255;
  ram[2829]  = 255;
  ram[2830]  = 255;
  ram[2831]  = 255;
  ram[2832]  = 236;
  ram[2833]  = 52;
  ram[2834]  = 0;
  ram[2835]  = 35;
  ram[2836]  = 208;
  ram[2837]  = 255;
  ram[2838]  = 35;
  ram[2839]  = 0;
  ram[2840]  = 208;
  ram[2841]  = 255;
  ram[2842]  = 255;
  ram[2843]  = 71;
  ram[2844]  = 0;
  ram[2845]  = 105;
  ram[2846]  = 137;
  ram[2847]  = 137;
  ram[2848]  = 137;
  ram[2849]  = 137;
  ram[2850]  = 137;
  ram[2851]  = 137;
  ram[2852]  = 137;
  ram[2853]  = 137;
  ram[2854]  = 0;
  ram[2855]  = 0;
  ram[2856]  = 255;
  ram[2857]  = 255;
  ram[2858]  = 255;
  ram[2859]  = 255;
  ram[2860]  = 255;
  ram[2861]  = 255;
  ram[2862]  = 255;
  ram[2863]  = 255;
  ram[2864]  = 255;
  ram[2865]  = 255;
  ram[2866]  = 255;
  ram[2867]  = 255;
  ram[2868]  = 255;
  ram[2869]  = 255;
  ram[2870]  = 255;
  ram[2871]  = 255;
  ram[2872]  = 255;
  ram[2873]  = 255;
  ram[2874]  = 255;
  ram[2875]  = 255;
  ram[2876]  = 255;
  ram[2877]  = 255;
  ram[2878]  = 255;
  ram[2879]  = 255;
  ram[2880]  = 255;
  ram[2881]  = 255;
  ram[2882]  = 255;
  ram[2883]  = 255;
  ram[2884]  = 255;
  ram[2885]  = 17;
  ram[2886]  = 0;
  ram[2887]  = 0;
  ram[2888]  = 221;
  ram[2889]  = 255;
  ram[2890]  = 255;
  ram[2891]  = 255;
  ram[2892]  = 255;
  ram[2893]  = 255;
  ram[2894]  = 255;
  ram[2895]  = 255;
  ram[2896]  = 255;
  ram[2897]  = 255;
  ram[2898]  = 255;
  ram[2899]  = 255;
  ram[2900]  = 255;
  ram[2901]  = 255;
  ram[2902]  = 255;
  ram[2903]  = 255;
  ram[2904]  = 255;
  ram[2905]  = 255;
  ram[2906]  = 255;
  ram[2907]  = 255;
  ram[2908]  = 255;
  ram[2909]  = 255;
  ram[2910]  = 255;
  ram[2911]  = 255;
  ram[2912]  = 255;
  ram[2913]  = 255;
  ram[2914]  = 255;
  ram[2915]  = 255;
  ram[2916]  = 255;
  ram[2917]  = 255;
  ram[2918]  = 255;
  ram[2919]  = 255;
  ram[2920]  = 255;
  ram[2921]  = 255;
  ram[2922]  = 255;
  ram[2923]  = 167;
  ram[2924]  = 0;
  ram[2925]  = 52;
  ram[2926]  = 255;
  ram[2927]  = 255;
  ram[2928]  = 255;
  ram[2929]  = 255;
  ram[2930]  = 255;
  ram[2931]  = 255;
  ram[2932]  = 255;
  ram[2933]  = 255;
  ram[2934]  = 71;
  ram[2935]  = 0;
  ram[2936]  = 137;
  ram[2937]  = 255;
  ram[2938]  = 255;
  ram[2939]  = 255;
  ram[2940]  = 255;
  ram[2941]  = 255;
  ram[2942]  = 255;
  ram[2943]  = 255;
  ram[2944]  = 255;
  ram[2945]  = 255;
  ram[2946]  = 255;
  ram[2947]  = 255;
  ram[2948]  = 255;
  ram[2949]  = 255;
  ram[2950]  = 255;
  ram[2951]  = 255;
  ram[2952]  = 255;
  ram[2953]  = 236;
  ram[2954]  = 71;
  ram[2955]  = 0;
  ram[2956]  = 17;
  ram[2957]  = 87;
  ram[2958]  = 0;
  ram[2959]  = 35;
  ram[2960]  = 255;
  ram[2961]  = 255;
  ram[2962]  = 255;
  ram[2963]  = 71;
  ram[2964]  = 0;
  ram[2965]  = 195;
  ram[2966]  = 255;
  ram[2967]  = 255;
  ram[2968]  = 255;
  ram[2969]  = 255;
  ram[2970]  = 255;
  ram[2971]  = 255;
  ram[2972]  = 255;
  ram[2973]  = 255;
  ram[2974]  = 0;
  ram[2975]  = 0;
  ram[2976]  = 255;
  ram[2977]  = 255;
  ram[2978]  = 255;
  ram[2979]  = 255;
  ram[2980]  = 255;
  ram[2981]  = 255;
  ram[2982]  = 255;
  ram[2983]  = 255;
  ram[2984]  = 255;
  ram[2985]  = 255;
  ram[2986]  = 255;
  ram[2987]  = 255;
  ram[2988]  = 255;
  ram[2989]  = 255;
  ram[2990]  = 255;
  ram[2991]  = 255;
  ram[2992]  = 255;
  ram[2993]  = 255;
  ram[2994]  = 255;
  ram[2995]  = 255;
  ram[2996]  = 255;
  ram[2997]  = 255;
  ram[2998]  = 255;
  ram[2999]  = 255;
  ram[3000]  = 255;
  ram[3001]  = 255;
  ram[3002]  = 255;
  ram[3003]  = 255;
  ram[3004]  = 255;
  ram[3005]  = 137;
  ram[3006]  = 0;
  ram[3007]  = 0;
  ram[3008]  = 52;
  ram[3009]  = 255;
  ram[3010]  = 255;
  ram[3011]  = 255;
  ram[3012]  = 255;
  ram[3013]  = 255;
  ram[3014]  = 255;
  ram[3015]  = 255;
  ram[3016]  = 255;
  ram[3017]  = 255;
  ram[3018]  = 255;
  ram[3019]  = 255;
  ram[3020]  = 255;
  ram[3021]  = 255;
  ram[3022]  = 255;
  ram[3023]  = 255;
  ram[3024]  = 255;
  ram[3025]  = 255;
  ram[3026]  = 255;
  ram[3027]  = 255;
  ram[3028]  = 255;
  ram[3029]  = 255;
  ram[3030]  = 255;
  ram[3031]  = 255;
  ram[3032]  = 255;
  ram[3033]  = 255;
  ram[3034]  = 255;
  ram[3035]  = 255;
  ram[3036]  = 255;
  ram[3037]  = 255;
  ram[3038]  = 255;
  ram[3039]  = 255;
  ram[3040]  = 255;
  ram[3041]  = 255;
  ram[3042]  = 255;
  ram[3043]  = 122;
  ram[3044]  = 0;
  ram[3045]  = 87;
  ram[3046]  = 255;
  ram[3047]  = 255;
  ram[3048]  = 255;
  ram[3049]  = 255;
  ram[3050]  = 255;
  ram[3051]  = 255;
  ram[3052]  = 255;
  ram[3053]  = 255;
  ram[3054]  = 71;
  ram[3055]  = 0;
  ram[3056]  = 137;
  ram[3057]  = 255;
  ram[3058]  = 255;
  ram[3059]  = 255;
  ram[3060]  = 255;
  ram[3061]  = 255;
  ram[3062]  = 255;
  ram[3063]  = 255;
  ram[3064]  = 255;
  ram[3065]  = 255;
  ram[3066]  = 255;
  ram[3067]  = 255;
  ram[3068]  = 255;
  ram[3069]  = 255;
  ram[3070]  = 255;
  ram[3071]  = 255;
  ram[3072]  = 255;
  ram[3073]  = 255;
  ram[3074]  = 255;
  ram[3075]  = 105;
  ram[3076]  = 0;
  ram[3077]  = 0;
  ram[3078]  = 0;
  ram[3079]  = 167;
  ram[3080]  = 255;
  ram[3081]  = 255;
  ram[3082]  = 255;
  ram[3083]  = 71;
  ram[3084]  = 0;
  ram[3085]  = 195;
  ram[3086]  = 255;
  ram[3087]  = 255;
  ram[3088]  = 255;
  ram[3089]  = 255;
  ram[3090]  = 255;
  ram[3091]  = 255;
  ram[3092]  = 255;
  ram[3093]  = 255;
  ram[3094]  = 0;
  ram[3095]  = 0;
  ram[3096]  = 255;
  ram[3097]  = 255;
  ram[3098]  = 255;
  ram[3099]  = 255;
  ram[3100]  = 255;
  ram[3101]  = 255;
  ram[3102]  = 255;
  ram[3103]  = 255;
  ram[3104]  = 255;
  ram[3105]  = 255;
  ram[3106]  = 255;
  ram[3107]  = 255;
  ram[3108]  = 255;
  ram[3109]  = 255;
  ram[3110]  = 255;
  ram[3111]  = 255;
  ram[3112]  = 255;
  ram[3113]  = 255;
  ram[3114]  = 255;
  ram[3115]  = 255;
  ram[3116]  = 255;
  ram[3117]  = 255;
  ram[3118]  = 255;
  ram[3119]  = 255;
  ram[3120]  = 255;
  ram[3121]  = 255;
  ram[3122]  = 255;
  ram[3123]  = 255;
  ram[3124]  = 255;
  ram[3125]  = 236;
  ram[3126]  = 35;
  ram[3127]  = 0;
  ram[3128]  = 0;
  ram[3129]  = 71;
  ram[3130]  = 236;
  ram[3131]  = 255;
  ram[3132]  = 255;
  ram[3133]  = 255;
  ram[3134]  = 255;
  ram[3135]  = 255;
  ram[3136]  = 255;
  ram[3137]  = 255;
  ram[3138]  = 255;
  ram[3139]  = 236;
  ram[3140]  = 255;
  ram[3141]  = 255;
  ram[3142]  = 255;
  ram[3143]  = 255;
  ram[3144]  = 255;
  ram[3145]  = 255;
  ram[3146]  = 255;
  ram[3147]  = 255;
  ram[3148]  = 255;
  ram[3149]  = 255;
  ram[3150]  = 255;
  ram[3151]  = 255;
  ram[3152]  = 255;
  ram[3153]  = 255;
  ram[3154]  = 255;
  ram[3155]  = 255;
  ram[3156]  = 255;
  ram[3157]  = 255;
  ram[3158]  = 255;
  ram[3159]  = 255;
  ram[3160]  = 255;
  ram[3161]  = 255;
  ram[3162]  = 255;
  ram[3163]  = 35;
  ram[3164]  = 0;
  ram[3165]  = 152;
  ram[3166]  = 255;
  ram[3167]  = 255;
  ram[3168]  = 255;
  ram[3169]  = 255;
  ram[3170]  = 255;
  ram[3171]  = 255;
  ram[3172]  = 255;
  ram[3173]  = 255;
  ram[3174]  = 71;
  ram[3175]  = 0;
  ram[3176]  = 137;
  ram[3177]  = 255;
  ram[3178]  = 255;
  ram[3179]  = 255;
  ram[3180]  = 255;
  ram[3181]  = 255;
  ram[3182]  = 255;
  ram[3183]  = 255;
  ram[3184]  = 255;
  ram[3185]  = 255;
  ram[3186]  = 255;
  ram[3187]  = 255;
  ram[3188]  = 255;
  ram[3189]  = 255;
  ram[3190]  = 255;
  ram[3191]  = 255;
  ram[3192]  = 255;
  ram[3193]  = 255;
  ram[3194]  = 255;
  ram[3195]  = 255;
  ram[3196]  = 71;
  ram[3197]  = 0;
  ram[3198]  = 0;
  ram[3199]  = 105;
  ram[3200]  = 255;
  ram[3201]  = 255;
  ram[3202]  = 255;
  ram[3203]  = 71;
  ram[3204]  = 0;
  ram[3205]  = 195;
  ram[3206]  = 255;
  ram[3207]  = 255;
  ram[3208]  = 255;
  ram[3209]  = 255;
  ram[3210]  = 255;
  ram[3211]  = 255;
  ram[3212]  = 255;
  ram[3213]  = 255;
  ram[3214]  = 0;
  ram[3215]  = 0;
  ram[3216]  = 255;
  ram[3217]  = 255;
  ram[3218]  = 255;
  ram[3219]  = 255;
  ram[3220]  = 255;
  ram[3221]  = 255;
  ram[3222]  = 255;
  ram[3223]  = 255;
  ram[3224]  = 255;
  ram[3225]  = 255;
  ram[3226]  = 255;
  ram[3227]  = 255;
  ram[3228]  = 255;
  ram[3229]  = 255;
  ram[3230]  = 255;
  ram[3231]  = 255;
  ram[3232]  = 255;
  ram[3233]  = 255;
  ram[3234]  = 255;
  ram[3235]  = 255;
  ram[3236]  = 255;
  ram[3237]  = 255;
  ram[3238]  = 255;
  ram[3239]  = 255;
  ram[3240]  = 255;
  ram[3241]  = 255;
  ram[3242]  = 255;
  ram[3243]  = 255;
  ram[3244]  = 255;
  ram[3245]  = 255;
  ram[3246]  = 208;
  ram[3247]  = 17;
  ram[3248]  = 0;
  ram[3249]  = 0;
  ram[3250]  = 17;
  ram[3251]  = 137;
  ram[3252]  = 208;
  ram[3253]  = 255;
  ram[3254]  = 255;
  ram[3255]  = 255;
  ram[3256]  = 195;
  ram[3257]  = 152;
  ram[3258]  = 52;
  ram[3259]  = 137;
  ram[3260]  = 255;
  ram[3261]  = 255;
  ram[3262]  = 255;
  ram[3263]  = 255;
  ram[3264]  = 255;
  ram[3265]  = 255;
  ram[3266]  = 255;
  ram[3267]  = 255;
  ram[3268]  = 255;
  ram[3269]  = 255;
  ram[3270]  = 255;
  ram[3271]  = 255;
  ram[3272]  = 255;
  ram[3273]  = 255;
  ram[3274]  = 255;
  ram[3275]  = 255;
  ram[3276]  = 255;
  ram[3277]  = 255;
  ram[3278]  = 255;
  ram[3279]  = 255;
  ram[3280]  = 255;
  ram[3281]  = 255;
  ram[3282]  = 167;
  ram[3283]  = 0;
  ram[3284]  = 0;
  ram[3285]  = 221;
  ram[3286]  = 255;
  ram[3287]  = 255;
  ram[3288]  = 255;
  ram[3289]  = 255;
  ram[3290]  = 255;
  ram[3291]  = 255;
  ram[3292]  = 255;
  ram[3293]  = 255;
  ram[3294]  = 71;
  ram[3295]  = 0;
  ram[3296]  = 137;
  ram[3297]  = 255;
  ram[3298]  = 255;
  ram[3299]  = 255;
  ram[3300]  = 255;
  ram[3301]  = 255;
  ram[3302]  = 255;
  ram[3303]  = 255;
  ram[3304]  = 255;
  ram[3305]  = 255;
  ram[3306]  = 255;
  ram[3307]  = 255;
  ram[3308]  = 255;
  ram[3309]  = 255;
  ram[3310]  = 255;
  ram[3311]  = 255;
  ram[3312]  = 255;
  ram[3313]  = 255;
  ram[3314]  = 255;
  ram[3315]  = 208;
  ram[3316]  = 0;
  ram[3317]  = 0;
  ram[3318]  = 0;
  ram[3319]  = 0;
  ram[3320]  = 105;
  ram[3321]  = 255;
  ram[3322]  = 255;
  ram[3323]  = 71;
  ram[3324]  = 0;
  ram[3325]  = 195;
  ram[3326]  = 255;
  ram[3327]  = 255;
  ram[3328]  = 255;
  ram[3329]  = 255;
  ram[3330]  = 255;
  ram[3331]  = 255;
  ram[3332]  = 255;
  ram[3333]  = 255;
  ram[3334]  = 0;
  ram[3335]  = 0;
  ram[3336]  = 255;
  ram[3337]  = 255;
  ram[3338]  = 255;
  ram[3339]  = 255;
  ram[3340]  = 255;
  ram[3341]  = 255;
  ram[3342]  = 255;
  ram[3343]  = 255;
  ram[3344]  = 255;
  ram[3345]  = 255;
  ram[3346]  = 255;
  ram[3347]  = 255;
  ram[3348]  = 255;
  ram[3349]  = 255;
  ram[3350]  = 255;
  ram[3351]  = 255;
  ram[3352]  = 255;
  ram[3353]  = 255;
  ram[3354]  = 255;
  ram[3355]  = 255;
  ram[3356]  = 255;
  ram[3357]  = 255;
  ram[3358]  = 255;
  ram[3359]  = 255;
  ram[3360]  = 255;
  ram[3361]  = 255;
  ram[3362]  = 255;
  ram[3363]  = 255;
  ram[3364]  = 255;
  ram[3365]  = 255;
  ram[3366]  = 255;
  ram[3367]  = 208;
  ram[3368]  = 52;
  ram[3369]  = 0;
  ram[3370]  = 0;
  ram[3371]  = 0;
  ram[3372]  = 0;
  ram[3373]  = 0;
  ram[3374]  = 0;
  ram[3375]  = 0;
  ram[3376]  = 0;
  ram[3377]  = 0;
  ram[3378]  = 0;
  ram[3379]  = 137;
  ram[3380]  = 255;
  ram[3381]  = 255;
  ram[3382]  = 255;
  ram[3383]  = 255;
  ram[3384]  = 255;
  ram[3385]  = 255;
  ram[3386]  = 255;
  ram[3387]  = 255;
  ram[3388]  = 255;
  ram[3389]  = 255;
  ram[3390]  = 255;
  ram[3391]  = 255;
  ram[3392]  = 255;
  ram[3393]  = 255;
  ram[3394]  = 255;
  ram[3395]  = 255;
  ram[3396]  = 255;
  ram[3397]  = 255;
  ram[3398]  = 255;
  ram[3399]  = 255;
  ram[3400]  = 255;
  ram[3401]  = 208;
  ram[3402]  = 17;
  ram[3403]  = 0;
  ram[3404]  = 105;
  ram[3405]  = 255;
  ram[3406]  = 255;
  ram[3407]  = 255;
  ram[3408]  = 255;
  ram[3409]  = 255;
  ram[3410]  = 255;
  ram[3411]  = 255;
  ram[3412]  = 255;
  ram[3413]  = 255;
  ram[3414]  = 71;
  ram[3415]  = 0;
  ram[3416]  = 137;
  ram[3417]  = 255;
  ram[3418]  = 255;
  ram[3419]  = 255;
  ram[3420]  = 255;
  ram[3421]  = 255;
  ram[3422]  = 255;
  ram[3423]  = 255;
  ram[3424]  = 255;
  ram[3425]  = 255;
  ram[3426]  = 255;
  ram[3427]  = 255;
  ram[3428]  = 255;
  ram[3429]  = 255;
  ram[3430]  = 255;
  ram[3431]  = 255;
  ram[3432]  = 255;
  ram[3433]  = 255;
  ram[3434]  = 236;
  ram[3435]  = 35;
  ram[3436]  = 0;
  ram[3437]  = 122;
  ram[3438]  = 167;
  ram[3439]  = 0;
  ram[3440]  = 0;
  ram[3441]  = 52;
  ram[3442]  = 236;
  ram[3443]  = 71;
  ram[3444]  = 0;
  ram[3445]  = 195;
  ram[3446]  = 255;
  ram[3447]  = 255;
  ram[3448]  = 255;
  ram[3449]  = 255;
  ram[3450]  = 255;
  ram[3451]  = 255;
  ram[3452]  = 255;
  ram[3453]  = 255;
  ram[3454]  = 0;
  ram[3455]  = 0;
  ram[3456]  = 255;
  ram[3457]  = 255;
  ram[3458]  = 255;
  ram[3459]  = 255;
  ram[3460]  = 255;
  ram[3461]  = 255;
  ram[3462]  = 255;
  ram[3463]  = 255;
  ram[3464]  = 255;
  ram[3465]  = 255;
  ram[3466]  = 255;
  ram[3467]  = 255;
  ram[3468]  = 255;
  ram[3469]  = 255;
  ram[3470]  = 255;
  ram[3471]  = 255;
  ram[3472]  = 255;
  ram[3473]  = 255;
  ram[3474]  = 255;
  ram[3475]  = 255;
  ram[3476]  = 255;
  ram[3477]  = 255;
  ram[3478]  = 255;
  ram[3479]  = 255;
  ram[3480]  = 255;
  ram[3481]  = 255;
  ram[3482]  = 255;
  ram[3483]  = 255;
  ram[3484]  = 255;
  ram[3485]  = 255;
  ram[3486]  = 255;
  ram[3487]  = 255;
  ram[3488]  = 255;
  ram[3489]  = 167;
  ram[3490]  = 52;
  ram[3491]  = 0;
  ram[3492]  = 0;
  ram[3493]  = 0;
  ram[3494]  = 0;
  ram[3495]  = 0;
  ram[3496]  = 0;
  ram[3497]  = 17;
  ram[3498]  = 105;
  ram[3499]  = 208;
  ram[3500]  = 255;
  ram[3501]  = 255;
  ram[3502]  = 255;
  ram[3503]  = 255;
  ram[3504]  = 255;
  ram[3505]  = 255;
  ram[3506]  = 255;
  ram[3507]  = 255;
  ram[3508]  = 255;
  ram[3509]  = 255;
  ram[3510]  = 255;
  ram[3511]  = 255;
  ram[3512]  = 255;
  ram[3513]  = 255;
  ram[3514]  = 255;
  ram[3515]  = 255;
  ram[3516]  = 255;
  ram[3517]  = 255;
  ram[3518]  = 255;
  ram[3519]  = 255;
  ram[3520]  = 208;
  ram[3521]  = 17;
  ram[3522]  = 0;
  ram[3523]  = 17;
  ram[3524]  = 236;
  ram[3525]  = 255;
  ram[3526]  = 255;
  ram[3527]  = 255;
  ram[3528]  = 255;
  ram[3529]  = 255;
  ram[3530]  = 255;
  ram[3531]  = 255;
  ram[3532]  = 255;
  ram[3533]  = 255;
  ram[3534]  = 71;
  ram[3535]  = 0;
  ram[3536]  = 137;
  ram[3537]  = 255;
  ram[3538]  = 255;
  ram[3539]  = 255;
  ram[3540]  = 255;
  ram[3541]  = 255;
  ram[3542]  = 255;
  ram[3543]  = 255;
  ram[3544]  = 255;
  ram[3545]  = 255;
  ram[3546]  = 255;
  ram[3547]  = 255;
  ram[3548]  = 255;
  ram[3549]  = 255;
  ram[3550]  = 255;
  ram[3551]  = 255;
  ram[3552]  = 255;
  ram[3553]  = 236;
  ram[3554]  = 52;
  ram[3555]  = 0;
  ram[3556]  = 52;
  ram[3557]  = 255;
  ram[3558]  = 255;
  ram[3559]  = 167;
  ram[3560]  = 0;
  ram[3561]  = 35;
  ram[3562]  = 236;
  ram[3563]  = 71;
  ram[3564]  = 0;
  ram[3565]  = 152;
  ram[3566]  = 195;
  ram[3567]  = 195;
  ram[3568]  = 195;
  ram[3569]  = 195;
  ram[3570]  = 195;
  ram[3571]  = 195;
  ram[3572]  = 195;
  ram[3573]  = 195;
  ram[3574]  = 0;
  ram[3575]  = 0;
  ram[3576]  = 255;
  ram[3577]  = 255;
  ram[3578]  = 255;
  ram[3579]  = 255;
  ram[3580]  = 255;
  ram[3581]  = 255;
  ram[3582]  = 255;
  ram[3583]  = 255;
  ram[3584]  = 255;
  ram[3585]  = 255;
  ram[3586]  = 255;
  ram[3587]  = 255;
  ram[3588]  = 255;
  ram[3589]  = 255;
  ram[3590]  = 255;
  ram[3591]  = 255;
  ram[3592]  = 255;
  ram[3593]  = 255;
  ram[3594]  = 255;
  ram[3595]  = 255;
  ram[3596]  = 255;
  ram[3597]  = 255;
  ram[3598]  = 255;
  ram[3599]  = 255;
  ram[3600]  = 255;
  ram[3601]  = 255;
  ram[3602]  = 255;
  ram[3603]  = 255;
  ram[3604]  = 255;
  ram[3605]  = 255;
  ram[3606]  = 255;
  ram[3607]  = 255;
  ram[3608]  = 255;
  ram[3609]  = 255;
  ram[3610]  = 255;
  ram[3611]  = 236;
  ram[3612]  = 195;
  ram[3613]  = 195;
  ram[3614]  = 195;
  ram[3615]  = 195;
  ram[3616]  = 208;
  ram[3617]  = 255;
  ram[3618]  = 255;
  ram[3619]  = 255;
  ram[3620]  = 255;
  ram[3621]  = 255;
  ram[3622]  = 255;
  ram[3623]  = 255;
  ram[3624]  = 255;
  ram[3625]  = 255;
  ram[3626]  = 255;
  ram[3627]  = 255;
  ram[3628]  = 255;
  ram[3629]  = 255;
  ram[3630]  = 255;
  ram[3631]  = 255;
  ram[3632]  = 255;
  ram[3633]  = 255;
  ram[3634]  = 255;
  ram[3635]  = 255;
  ram[3636]  = 255;
  ram[3637]  = 255;
  ram[3638]  = 255;
  ram[3639]  = 137;
  ram[3640]  = 0;
  ram[3641]  = 0;
  ram[3642]  = 17;
  ram[3643]  = 208;
  ram[3644]  = 255;
  ram[3645]  = 255;
  ram[3646]  = 255;
  ram[3647]  = 255;
  ram[3648]  = 255;
  ram[3649]  = 255;
  ram[3650]  = 255;
  ram[3651]  = 255;
  ram[3652]  = 255;
  ram[3653]  = 255;
  ram[3654]  = 71;
  ram[3655]  = 0;
  ram[3656]  = 137;
  ram[3657]  = 255;
  ram[3658]  = 255;
  ram[3659]  = 255;
  ram[3660]  = 255;
  ram[3661]  = 255;
  ram[3662]  = 255;
  ram[3663]  = 255;
  ram[3664]  = 255;
  ram[3665]  = 255;
  ram[3666]  = 255;
  ram[3667]  = 255;
  ram[3668]  = 255;
  ram[3669]  = 255;
  ram[3670]  = 255;
  ram[3671]  = 255;
  ram[3672]  = 208;
  ram[3673]  = 52;
  ram[3674]  = 0;
  ram[3675]  = 52;
  ram[3676]  = 236;
  ram[3677]  = 255;
  ram[3678]  = 255;
  ram[3679]  = 255;
  ram[3680]  = 167;
  ram[3681]  = 208;
  ram[3682]  = 255;
  ram[3683]  = 71;
  ram[3684]  = 0;
  ram[3685]  = 0;
  ram[3686]  = 0;
  ram[3687]  = 0;
  ram[3688]  = 0;
  ram[3689]  = 0;
  ram[3690]  = 0;
  ram[3691]  = 0;
  ram[3692]  = 0;
  ram[3693]  = 0;
  ram[3694]  = 0;
  ram[3695]  = 0;
  ram[3696]  = 255;
  ram[3697]  = 255;
  ram[3698]  = 255;
  ram[3699]  = 255;
  ram[3700]  = 255;
  ram[3701]  = 255;
  ram[3702]  = 255;
  ram[3703]  = 255;
  ram[3704]  = 255;
  ram[3705]  = 255;
  ram[3706]  = 255;
  ram[3707]  = 255;
  ram[3708]  = 255;
  ram[3709]  = 255;
  ram[3710]  = 255;
  ram[3711]  = 255;
  ram[3712]  = 255;
  ram[3713]  = 255;
  ram[3714]  = 255;
  ram[3715]  = 255;
  ram[3716]  = 255;
  ram[3717]  = 255;
  ram[3718]  = 255;
  ram[3719]  = 255;
  ram[3720]  = 255;
  ram[3721]  = 255;
  ram[3722]  = 255;
  ram[3723]  = 255;
  ram[3724]  = 255;
  ram[3725]  = 255;
  ram[3726]  = 255;
  ram[3727]  = 255;
  ram[3728]  = 255;
  ram[3729]  = 255;
  ram[3730]  = 255;
  ram[3731]  = 255;
  ram[3732]  = 255;
  ram[3733]  = 255;
  ram[3734]  = 255;
  ram[3735]  = 255;
  ram[3736]  = 255;
  ram[3737]  = 255;
  ram[3738]  = 255;
  ram[3739]  = 255;
  ram[3740]  = 255;
  ram[3741]  = 255;
  ram[3742]  = 255;
  ram[3743]  = 255;
  ram[3744]  = 255;
  ram[3745]  = 255;
  ram[3746]  = 255;
  ram[3747]  = 255;
  ram[3748]  = 255;
  ram[3749]  = 255;
  ram[3750]  = 255;
  ram[3751]  = 255;
  ram[3752]  = 255;
  ram[3753]  = 255;
  ram[3754]  = 255;
  ram[3755]  = 255;
  ram[3756]  = 255;
  ram[3757]  = 195;
  ram[3758]  = 35;
  ram[3759]  = 0;
  ram[3760]  = 0;
  ram[3761]  = 52;
  ram[3762]  = 208;
  ram[3763]  = 255;
  ram[3764]  = 255;
  ram[3765]  = 255;
  ram[3766]  = 255;
  ram[3767]  = 255;
  ram[3768]  = 255;
  ram[3769]  = 255;
  ram[3770]  = 255;
  ram[3771]  = 255;
  ram[3772]  = 255;
  ram[3773]  = 255;
  ram[3774]  = 71;
  ram[3775]  = 0;
  ram[3776]  = 137;
  ram[3777]  = 255;
  ram[3778]  = 255;
  ram[3779]  = 255;
  ram[3780]  = 255;
  ram[3781]  = 255;
  ram[3782]  = 255;
  ram[3783]  = 255;
  ram[3784]  = 255;
  ram[3785]  = 255;
  ram[3786]  = 255;
  ram[3787]  = 255;
  ram[3788]  = 255;
  ram[3789]  = 255;
  ram[3790]  = 255;
  ram[3791]  = 221;
  ram[3792]  = 17;
  ram[3793]  = 0;
  ram[3794]  = 52;
  ram[3795]  = 236;
  ram[3796]  = 255;
  ram[3797]  = 255;
  ram[3798]  = 255;
  ram[3799]  = 255;
  ram[3800]  = 255;
  ram[3801]  = 255;
  ram[3802]  = 255;
  ram[3803]  = 71;
  ram[3804]  = 0;
  ram[3805]  = 52;
  ram[3806]  = 71;
  ram[3807]  = 71;
  ram[3808]  = 71;
  ram[3809]  = 71;
  ram[3810]  = 71;
  ram[3811]  = 71;
  ram[3812]  = 71;
  ram[3813]  = 71;
  ram[3814]  = 0;
  ram[3815]  = 0;
  ram[3816]  = 255;
  ram[3817]  = 255;
  ram[3818]  = 255;
  ram[3819]  = 255;
  ram[3820]  = 255;
  ram[3821]  = 255;
  ram[3822]  = 255;
  ram[3823]  = 255;
  ram[3824]  = 255;
  ram[3825]  = 255;
  ram[3826]  = 255;
  ram[3827]  = 255;
  ram[3828]  = 255;
  ram[3829]  = 255;
  ram[3830]  = 255;
  ram[3831]  = 255;
  ram[3832]  = 255;
  ram[3833]  = 255;
  ram[3834]  = 255;
  ram[3835]  = 255;
  ram[3836]  = 255;
  ram[3837]  = 255;
  ram[3838]  = 255;
  ram[3839]  = 255;
  ram[3840]  = 255;
  ram[3841]  = 255;
  ram[3842]  = 255;
  ram[3843]  = 255;
  ram[3844]  = 255;
  ram[3845]  = 255;
  ram[3846]  = 255;
  ram[3847]  = 255;
  ram[3848]  = 255;
  ram[3849]  = 255;
  ram[3850]  = 255;
  ram[3851]  = 255;
  ram[3852]  = 255;
  ram[3853]  = 255;
  ram[3854]  = 255;
  ram[3855]  = 255;
  ram[3856]  = 255;
  ram[3857]  = 255;
  ram[3858]  = 255;
  ram[3859]  = 255;
  ram[3860]  = 255;
  ram[3861]  = 255;
  ram[3862]  = 255;
  ram[3863]  = 255;
  ram[3864]  = 255;
  ram[3865]  = 255;
  ram[3866]  = 255;
  ram[3867]  = 255;
  ram[3868]  = 255;
  ram[3869]  = 255;
  ram[3870]  = 255;
  ram[3871]  = 255;
  ram[3872]  = 255;
  ram[3873]  = 255;
  ram[3874]  = 255;
  ram[3875]  = 255;
  ram[3876]  = 255;
  ram[3877]  = 208;
  ram[3878]  = 17;
  ram[3879]  = 0;
  ram[3880]  = 122;
  ram[3881]  = 236;
  ram[3882]  = 255;
  ram[3883]  = 255;
  ram[3884]  = 255;
  ram[3885]  = 255;
  ram[3886]  = 255;
  ram[3887]  = 255;
  ram[3888]  = 255;
  ram[3889]  = 255;
  ram[3890]  = 255;
  ram[3891]  = 255;
  ram[3892]  = 255;
  ram[3893]  = 255;
  ram[3894]  = 71;
  ram[3895]  = 0;
  ram[3896]  = 137;
  ram[3897]  = 255;
  ram[3898]  = 255;
  ram[3899]  = 255;
  ram[3900]  = 255;
  ram[3901]  = 255;
  ram[3902]  = 255;
  ram[3903]  = 255;
  ram[3904]  = 255;
  ram[3905]  = 255;
  ram[3906]  = 255;
  ram[3907]  = 255;
  ram[3908]  = 255;
  ram[3909]  = 255;
  ram[3910]  = 255;
  ram[3911]  = 255;
  ram[3912]  = 87;
  ram[3913]  = 71;
  ram[3914]  = 236;
  ram[3915]  = 255;
  ram[3916]  = 255;
  ram[3917]  = 255;
  ram[3918]  = 255;
  ram[3919]  = 255;
  ram[3920]  = 255;
  ram[3921]  = 255;
  ram[3922]  = 255;
  ram[3923]  = 71;
  ram[3924]  = 0;
  ram[3925]  = 195;
  ram[3926]  = 255;
  ram[3927]  = 255;
  ram[3928]  = 255;
  ram[3929]  = 255;
  ram[3930]  = 255;
  ram[3931]  = 255;
  ram[3932]  = 255;
  ram[3933]  = 255;
  ram[3934]  = 0;
  ram[3935]  = 0;
  ram[3936]  = 255;
  ram[3937]  = 255;
  ram[3938]  = 255;
  ram[3939]  = 255;
  ram[3940]  = 255;
  ram[3941]  = 255;
  ram[3942]  = 255;
  ram[3943]  = 255;
  ram[3944]  = 255;
  ram[3945]  = 255;
  ram[3946]  = 255;
  ram[3947]  = 255;
  ram[3948]  = 255;
  ram[3949]  = 255;
  ram[3950]  = 255;
  ram[3951]  = 255;
  ram[3952]  = 255;
  ram[3953]  = 255;
  ram[3954]  = 255;
  ram[3955]  = 255;
  ram[3956]  = 255;
  ram[3957]  = 255;
  ram[3958]  = 255;
  ram[3959]  = 255;
  ram[3960]  = 255;
  ram[3961]  = 255;
  ram[3962]  = 255;
  ram[3963]  = 255;
  ram[3964]  = 255;
  ram[3965]  = 255;
  ram[3966]  = 255;
  ram[3967]  = 255;
  ram[3968]  = 255;
  ram[3969]  = 255;
  ram[3970]  = 255;
  ram[3971]  = 255;
  ram[3972]  = 255;
  ram[3973]  = 255;
  ram[3974]  = 255;
  ram[3975]  = 255;
  ram[3976]  = 255;
  ram[3977]  = 255;
  ram[3978]  = 255;
  ram[3979]  = 255;
  ram[3980]  = 255;
  ram[3981]  = 255;
  ram[3982]  = 255;
  ram[3983]  = 255;
  ram[3984]  = 255;
  ram[3985]  = 255;
  ram[3986]  = 255;
  ram[3987]  = 255;
  ram[3988]  = 255;
  ram[3989]  = 255;
  ram[3990]  = 255;
  ram[3991]  = 255;
  ram[3992]  = 255;
  ram[3993]  = 255;
  ram[3994]  = 255;
  ram[3995]  = 255;
  ram[3996]  = 255;
  ram[3997]  = 255;
  ram[3998]  = 181;
  ram[3999]  = 195;
  ram[4000]  = 255;
  ram[4001]  = 255;
  ram[4002]  = 255;
  ram[4003]  = 255;
  ram[4004]  = 255;
  ram[4005]  = 255;
  ram[4006]  = 255;
  ram[4007]  = 255;
  ram[4008]  = 255;
  ram[4009]  = 255;
  ram[4010]  = 255;
  ram[4011]  = 255;
  ram[4012]  = 255;
  ram[4013]  = 255;
  ram[4014]  = 208;
  ram[4015]  = 195;
  ram[4016]  = 221;
  ram[4017]  = 255;
  ram[4018]  = 255;
  ram[4019]  = 255;
  ram[4020]  = 255;
  ram[4021]  = 255;
  ram[4022]  = 255;
  ram[4023]  = 255;
  ram[4024]  = 255;
  ram[4025]  = 255;
  ram[4026]  = 255;
  ram[4027]  = 255;
  ram[4028]  = 255;
  ram[4029]  = 255;
  ram[4030]  = 255;
  ram[4031]  = 255;
  ram[4032]  = 236;
  ram[4033]  = 255;
  ram[4034]  = 255;
  ram[4035]  = 255;
  ram[4036]  = 255;
  ram[4037]  = 255;
  ram[4038]  = 255;
  ram[4039]  = 255;
  ram[4040]  = 255;
  ram[4041]  = 255;
  ram[4042]  = 255;
  ram[4043]  = 167;
  ram[4044]  = 137;
  ram[4045]  = 221;
  ram[4046]  = 255;
  ram[4047]  = 255;
  ram[4048]  = 255;
  ram[4049]  = 255;
  ram[4050]  = 255;
  ram[4051]  = 255;
  ram[4052]  = 255;
  ram[4053]  = 255;
  ram[4054]  = 137;
  ram[4055]  = 137;
  ram[4056]  = 255;
  ram[4057]  = 255;
  ram[4058]  = 255;
  ram[4059]  = 255;
  ram[4060]  = 255;
  ram[4061]  = 255;
  ram[4062]  = 255;
  ram[4063]  = 255;
  ram[4064]  = 255;
  ram[4065]  = 255;
  ram[4066]  = 255;
  ram[4067]  = 255;
  ram[4068]  = 255;
  ram[4069]  = 255;
  ram[4070]  = 255;
  ram[4071]  = 255;
  ram[4072]  = 255;
  ram[4073]  = 255;
  ram[4074]  = 255;
  ram[4075]  = 255;
  ram[4076]  = 255;
  ram[4077]  = 255;
  ram[4078]  = 255;
  ram[4079]  = 255;
  ram[4080]  = 255;
  ram[4081]  = 255;
  ram[4082]  = 255;
  ram[4083]  = 255;
  ram[4084]  = 255;
  ram[4085]  = 255;
  ram[4086]  = 255;
  ram[4087]  = 255;
  ram[4088]  = 255;
  ram[4089]  = 255;
  ram[4090]  = 255;
  ram[4091]  = 255;
  ram[4092]  = 255;
  ram[4093]  = 255;
  ram[4094]  = 255;
  ram[4095]  = 255;
  ram[4096]  = 255;
  ram[4097]  = 255;
  ram[4098]  = 255;
  ram[4099]  = 255;
  ram[4100]  = 255;
  ram[4101]  = 255;
  ram[4102]  = 255;
  ram[4103]  = 255;
  ram[4104]  = 255;
  ram[4105]  = 255;
  ram[4106]  = 255;
  ram[4107]  = 255;
  ram[4108]  = 255;
  ram[4109]  = 255;
  ram[4110]  = 255;
  ram[4111]  = 255;
  ram[4112]  = 255;
  ram[4113]  = 255;
  ram[4114]  = 255;
  ram[4115]  = 255;
  ram[4116]  = 255;
  ram[4117]  = 255;
  ram[4118]  = 255;
  ram[4119]  = 255;
  ram[4120]  = 255;
  ram[4121]  = 255;
  ram[4122]  = 255;
  ram[4123]  = 255;
  ram[4124]  = 255;
  ram[4125]  = 255;
  ram[4126]  = 255;
  ram[4127]  = 255;
  ram[4128]  = 255;
  ram[4129]  = 255;
  ram[4130]  = 255;
  ram[4131]  = 255;
  ram[4132]  = 255;
  ram[4133]  = 255;
  ram[4134]  = 255;
  ram[4135]  = 255;
  ram[4136]  = 255;
  ram[4137]  = 255;
  ram[4138]  = 255;
  ram[4139]  = 255;
  ram[4140]  = 255;
  ram[4141]  = 255;
  ram[4142]  = 255;
  ram[4143]  = 255;
  ram[4144]  = 255;
  ram[4145]  = 255;
  ram[4146]  = 255;
  ram[4147]  = 255;
  ram[4148]  = 255;
  ram[4149]  = 255;
  ram[4150]  = 255;
  ram[4151]  = 255;
  ram[4152]  = 255;
  ram[4153]  = 255;
  ram[4154]  = 255;
  ram[4155]  = 255;
  ram[4156]  = 255;
  ram[4157]  = 255;
  ram[4158]  = 255;
  ram[4159]  = 255;
  ram[4160]  = 255;
  ram[4161]  = 255;
  ram[4162]  = 255;
  ram[4163]  = 255;
  ram[4164]  = 255;
  ram[4165]  = 255;
  ram[4166]  = 255;
  ram[4167]  = 255;
  ram[4168]  = 255;
  ram[4169]  = 255;
  ram[4170]  = 255;
  ram[4171]  = 255;
  ram[4172]  = 255;
  ram[4173]  = 255;
  ram[4174]  = 255;
  ram[4175]  = 255;
  ram[4176]  = 255;
  ram[4177]  = 255;
  ram[4178]  = 255;
  ram[4179]  = 255;
  ram[4180]  = 255;
  ram[4181]  = 255;
  ram[4182]  = 255;
  ram[4183]  = 255;
  ram[4184]  = 255;
  ram[4185]  = 255;
  ram[4186]  = 255;
  ram[4187]  = 255;
  ram[4188]  = 255;
  ram[4189]  = 255;
  ram[4190]  = 255;
  ram[4191]  = 255;
  ram[4192]  = 255;
  ram[4193]  = 255;
  ram[4194]  = 255;
  ram[4195]  = 255;
  ram[4196]  = 255;
  ram[4197]  = 255;
  ram[4198]  = 255;
  ram[4199]  = 255;
  ram[4200]  = 255;
  ram[4201]  = 255;
  ram[4202]  = 255;
  ram[4203]  = 255;
  ram[4204]  = 255;
  ram[4205]  = 255;
  ram[4206]  = 255;
  ram[4207]  = 255;
  ram[4208]  = 255;
  ram[4209]  = 255;
  ram[4210]  = 255;
  ram[4211]  = 255;
  ram[4212]  = 255;
  ram[4213]  = 255;
  ram[4214]  = 255;
  ram[4215]  = 255;
  ram[4216]  = 255;
  ram[4217]  = 255;
  ram[4218]  = 255;
  ram[4219]  = 255;
  ram[4220]  = 255;
  ram[4221]  = 255;
  ram[4222]  = 255;
  ram[4223]  = 255;
  ram[4224]  = 255;
  ram[4225]  = 255;
  ram[4226]  = 255;
  ram[4227]  = 255;
  ram[4228]  = 255;
  ram[4229]  = 255;
  ram[4230]  = 255;
  ram[4231]  = 255;
  ram[4232]  = 255;
  ram[4233]  = 255;
  ram[4234]  = 255;
  ram[4235]  = 255;
  ram[4236]  = 255;
  ram[4237]  = 255;
  ram[4238]  = 255;
  ram[4239]  = 255;
  ram[4240]  = 255;
  ram[4241]  = 255;
  ram[4242]  = 255;
  ram[4243]  = 255;
  ram[4244]  = 255;
  ram[4245]  = 255;
  ram[4246]  = 255;
  ram[4247]  = 255;
  ram[4248]  = 255;
  ram[4249]  = 255;
  ram[4250]  = 255;
  ram[4251]  = 255;
  ram[4252]  = 255;
  ram[4253]  = 255;
  ram[4254]  = 255;
  ram[4255]  = 255;
  ram[4256]  = 255;
  ram[4257]  = 255;
  ram[4258]  = 255;
  ram[4259]  = 255;
  ram[4260]  = 255;
  ram[4261]  = 255;
  ram[4262]  = 255;
  ram[4263]  = 255;
  ram[4264]  = 255;
  ram[4265]  = 255;
  ram[4266]  = 255;
  ram[4267]  = 255;
  ram[4268]  = 255;
  ram[4269]  = 255;
  ram[4270]  = 255;
  ram[4271]  = 255;
  ram[4272]  = 255;
  ram[4273]  = 255;
  ram[4274]  = 255;
  ram[4275]  = 255;
  ram[4276]  = 255;
  ram[4277]  = 255;
  ram[4278]  = 255;
  ram[4279]  = 255;
  ram[4280]  = 255;
  ram[4281]  = 255;
  ram[4282]  = 255;
  ram[4283]  = 255;
  ram[4284]  = 255;
  ram[4285]  = 255;
  ram[4286]  = 255;
  ram[4287]  = 255;
  ram[4288]  = 255;
  ram[4289]  = 255;
  ram[4290]  = 255;
  ram[4291]  = 255;
  ram[4292]  = 255;
  ram[4293]  = 255;
  ram[4294]  = 255;
  ram[4295]  = 255;
  ram[4296]  = 255;
  ram[4297]  = 255;
  ram[4298]  = 255;
  ram[4299]  = 255;
  ram[4300]  = 255;
  ram[4301]  = 255;
  ram[4302]  = 255;
  ram[4303]  = 255;
  ram[4304]  = 255;
  ram[4305]  = 255;
  ram[4306]  = 255;
  ram[4307]  = 255;
  ram[4308]  = 255;
  ram[4309]  = 255;
  ram[4310]  = 255;
  ram[4311]  = 255;
  ram[4312]  = 255;
  ram[4313]  = 255;
  ram[4314]  = 255;
  ram[4315]  = 255;
  ram[4316]  = 255;
  ram[4317]  = 255;
  ram[4318]  = 255;
  ram[4319]  = 255;
  ram[4320]  = 255;
  ram[4321]  = 255;
  ram[4322]  = 255;
  ram[4323]  = 255;
  ram[4324]  = 255;
  ram[4325]  = 255;
  ram[4326]  = 255;
  ram[4327]  = 255;
  ram[4328]  = 255;
  ram[4329]  = 255;
  ram[4330]  = 255;
  ram[4331]  = 255;
  ram[4332]  = 255;
  ram[4333]  = 255;
  ram[4334]  = 255;
  ram[4335]  = 255;
  ram[4336]  = 255;
  ram[4337]  = 255;
  ram[4338]  = 255;
  ram[4339]  = 255;
  ram[4340]  = 255;
  ram[4341]  = 255;
  ram[4342]  = 255;
  ram[4343]  = 255;
  ram[4344]  = 255;
  ram[4345]  = 255;
  ram[4346]  = 255;
  ram[4347]  = 255;
  ram[4348]  = 255;
  ram[4349]  = 255;
  ram[4350]  = 255;
  ram[4351]  = 255;
  ram[4352]  = 255;
  ram[4353]  = 255;
  ram[4354]  = 255;
  ram[4355]  = 255;
  ram[4356]  = 255;
  ram[4357]  = 255;
  ram[4358]  = 255;
  ram[4359]  = 255;
  ram[4360]  = 255;
  ram[4361]  = 255;
  ram[4362]  = 255;
  ram[4363]  = 255;
  ram[4364]  = 255;
  ram[4365]  = 255;
  ram[4366]  = 255;
  ram[4367]  = 255;
  ram[4368]  = 255;
  ram[4369]  = 255;
  ram[4370]  = 255;
  ram[4371]  = 255;
  ram[4372]  = 255;
  ram[4373]  = 255;
  ram[4374]  = 255;
  ram[4375]  = 255;
  ram[4376]  = 255;
  ram[4377]  = 255;
  ram[4378]  = 255;
  ram[4379]  = 255;
  ram[4380]  = 255;
  ram[4381]  = 255;
  ram[4382]  = 255;
  ram[4383]  = 255;
  ram[4384]  = 255;
  ram[4385]  = 255;
  ram[4386]  = 255;
  ram[4387]  = 255;
  ram[4388]  = 255;
  ram[4389]  = 255;
  ram[4390]  = 255;
  ram[4391]  = 255;
  ram[4392]  = 255;
  ram[4393]  = 255;
  ram[4394]  = 255;
  ram[4395]  = 255;
  ram[4396]  = 255;
  ram[4397]  = 255;
  ram[4398]  = 255;
  ram[4399]  = 255;
  ram[4400]  = 255;
  ram[4401]  = 255;
  ram[4402]  = 255;
  ram[4403]  = 255;
  ram[4404]  = 255;
  ram[4405]  = 255;
  ram[4406]  = 255;
  ram[4407]  = 255;
  ram[4408]  = 255;
  ram[4409]  = 255;
  ram[4410]  = 255;
  ram[4411]  = 255;
  ram[4412]  = 255;
  ram[4413]  = 255;
  ram[4414]  = 255;
  ram[4415]  = 255;
  ram[4416]  = 255;
  ram[4417]  = 255;
  ram[4418]  = 255;
  ram[4419]  = 255;
  ram[4420]  = 255;
  ram[4421]  = 255;
  ram[4422]  = 255;
  ram[4423]  = 255;
  ram[4424]  = 255;
  ram[4425]  = 255;
  ram[4426]  = 255;
  ram[4427]  = 255;
  ram[4428]  = 255;
  ram[4429]  = 255;
  ram[4430]  = 255;
  ram[4431]  = 255;
  ram[4432]  = 255;
  ram[4433]  = 255;
  ram[4434]  = 255;
  ram[4435]  = 255;
  ram[4436]  = 255;
  ram[4437]  = 255;
  ram[4438]  = 255;
  ram[4439]  = 255;
  ram[4440]  = 255;
  ram[4441]  = 255;
  ram[4442]  = 255;
  ram[4443]  = 255;
  ram[4444]  = 255;
  ram[4445]  = 255;
  ram[4446]  = 255;
  ram[4447]  = 255;
  ram[4448]  = 255;
  ram[4449]  = 255;
  ram[4450]  = 255;
  ram[4451]  = 255;
  ram[4452]  = 255;
  ram[4453]  = 255;
  ram[4454]  = 255;
  ram[4455]  = 255;
  ram[4456]  = 255;
  ram[4457]  = 255;
  ram[4458]  = 255;
  ram[4459]  = 255;
  ram[4460]  = 255;
  ram[4461]  = 255;
  ram[4462]  = 255;
  ram[4463]  = 255;
  ram[4464]  = 255;
  ram[4465]  = 255;
  ram[4466]  = 255;
  ram[4467]  = 255;
  ram[4468]  = 255;
  ram[4469]  = 255;
  ram[4470]  = 255;
  ram[4471]  = 255;
  ram[4472]  = 255;
  ram[4473]  = 255;
  ram[4474]  = 255;
  ram[4475]  = 255;
  ram[4476]  = 255;
  ram[4477]  = 255;
  ram[4478]  = 255;
  ram[4479]  = 255;
  ram[4480]  = 255;
  ram[4481]  = 255;
  ram[4482]  = 255;
  ram[4483]  = 255;
  ram[4484]  = 255;
  ram[4485]  = 255;
  ram[4486]  = 255;
  ram[4487]  = 255;
  ram[4488]  = 255;
  ram[4489]  = 255;
  ram[4490]  = 255;
  ram[4491]  = 255;
  ram[4492]  = 255;
  ram[4493]  = 255;
  ram[4494]  = 255;
  ram[4495]  = 255;
  ram[4496]  = 255;
  ram[4497]  = 255;
  ram[4498]  = 255;
  ram[4499]  = 255;
  ram[4500]  = 255;
  ram[4501]  = 255;
  ram[4502]  = 255;
  ram[4503]  = 255;
  ram[4504]  = 255;
  ram[4505]  = 255;
  ram[4506]  = 255;
  ram[4507]  = 255;
  ram[4508]  = 255;
  ram[4509]  = 255;
  ram[4510]  = 255;
  ram[4511]  = 255;
  ram[4512]  = 255;
  ram[4513]  = 255;
  ram[4514]  = 255;
  ram[4515]  = 255;
  ram[4516]  = 255;
  ram[4517]  = 255;
  ram[4518]  = 255;
  ram[4519]  = 255;
  ram[4520]  = 255;
  ram[4521]  = 255;
  ram[4522]  = 255;
  ram[4523]  = 255;
  ram[4524]  = 255;
  ram[4525]  = 255;
  ram[4526]  = 255;
  ram[4527]  = 255;
  ram[4528]  = 255;
  ram[4529]  = 255;
  ram[4530]  = 255;
  ram[4531]  = 255;
  ram[4532]  = 255;
  ram[4533]  = 255;
  ram[4534]  = 255;
  ram[4535]  = 255;
  ram[4536]  = 255;
  ram[4537]  = 255;
  ram[4538]  = 255;
  ram[4539]  = 255;
  ram[4540]  = 255;
  ram[4541]  = 255;
  ram[4542]  = 255;
  ram[4543]  = 255;
  ram[4544]  = 255;
  ram[4545]  = 255;
  ram[4546]  = 255;
  ram[4547]  = 255;
  ram[4548]  = 255;
  ram[4549]  = 255;
  ram[4550]  = 255;
  ram[4551]  = 255;
  ram[4552]  = 255;
  ram[4553]  = 255;
  ram[4554]  = 255;
  ram[4555]  = 255;
  ram[4556]  = 255;
  ram[4557]  = 255;
  ram[4558]  = 255;
  ram[4559]  = 255;
  ram[4560]  = 255;
  ram[4561]  = 255;
  ram[4562]  = 255;
  ram[4563]  = 255;
  ram[4564]  = 255;
  ram[4565]  = 255;
  ram[4566]  = 255;
  ram[4567]  = 255;
  ram[4568]  = 255;
  ram[4569]  = 255;
  ram[4570]  = 255;
  ram[4571]  = 255;
  ram[4572]  = 255;
  ram[4573]  = 255;
  ram[4574]  = 255;
  ram[4575]  = 255;
  ram[4576]  = 255;
  ram[4577]  = 255;
  ram[4578]  = 255;
  ram[4579]  = 255;
  ram[4580]  = 255;
  ram[4581]  = 255;
  ram[4582]  = 255;
  ram[4583]  = 255;
  ram[4584]  = 255;
  ram[4585]  = 255;
  ram[4586]  = 255;
  ram[4587]  = 255;
  ram[4588]  = 255;
  ram[4589]  = 255;
  ram[4590]  = 255;
  ram[4591]  = 255;
  ram[4592]  = 255;
  ram[4593]  = 255;
  ram[4594]  = 255;
  ram[4595]  = 255;
  ram[4596]  = 255;
  ram[4597]  = 255;
  ram[4598]  = 255;
  ram[4599]  = 255;
  ram[4600]  = 255;
  ram[4601]  = 255;
  ram[4602]  = 255;
  ram[4603]  = 255;
  ram[4604]  = 255;
  ram[4605]  = 255;
  ram[4606]  = 255;
  ram[4607]  = 255;
  ram[4608]  = 255;
  ram[4609]  = 255;
  ram[4610]  = 255;
  ram[4611]  = 255;
  ram[4612]  = 255;
  ram[4613]  = 255;
  ram[4614]  = 255;
  ram[4615]  = 255;
  ram[4616]  = 255;
  ram[4617]  = 255;
  ram[4618]  = 255;
  ram[4619]  = 255;
  ram[4620]  = 255;
  ram[4621]  = 255;
  ram[4622]  = 255;
  ram[4623]  = 255;
  ram[4624]  = 255;
  ram[4625]  = 255;
  ram[4626]  = 255;
  ram[4627]  = 255;
  ram[4628]  = 255;
  ram[4629]  = 255;
  ram[4630]  = 255;
  ram[4631]  = 255;
  ram[4632]  = 255;
  ram[4633]  = 255;
  ram[4634]  = 255;
  ram[4635]  = 255;
  ram[4636]  = 255;
  ram[4637]  = 255;
  ram[4638]  = 255;
  ram[4639]  = 255;
  ram[4640]  = 255;
  ram[4641]  = 255;
  ram[4642]  = 255;
  ram[4643]  = 255;
  ram[4644]  = 255;
  ram[4645]  = 255;
  ram[4646]  = 255;
  ram[4647]  = 255;
  ram[4648]  = 255;
  ram[4649]  = 255;
  ram[4650]  = 255;
  ram[4651]  = 255;
  ram[4652]  = 255;
  ram[4653]  = 255;
  ram[4654]  = 255;
  ram[4655]  = 255;
  ram[4656]  = 255;
  ram[4657]  = 255;
  ram[4658]  = 255;
  ram[4659]  = 255;
  ram[4660]  = 255;
  ram[4661]  = 255;
  ram[4662]  = 255;
  ram[4663]  = 255;
  ram[4664]  = 255;
  ram[4665]  = 255;
  ram[4666]  = 255;
  ram[4667]  = 255;
  ram[4668]  = 255;
  ram[4669]  = 255;
  ram[4670]  = 255;
  ram[4671]  = 255;
  ram[4672]  = 255;
  ram[4673]  = 255;
  ram[4674]  = 255;
  ram[4675]  = 255;
  ram[4676]  = 255;
  ram[4677]  = 255;
  ram[4678]  = 255;
  ram[4679]  = 255;
  ram[4680]  = 255;
  ram[4681]  = 255;
  ram[4682]  = 255;
  ram[4683]  = 255;
  ram[4684]  = 255;
  ram[4685]  = 255;
  ram[4686]  = 255;
  ram[4687]  = 255;
  ram[4688]  = 255;
  ram[4689]  = 255;
  ram[4690]  = 255;
  ram[4691]  = 255;
  ram[4692]  = 255;
  ram[4693]  = 255;
  ram[4694]  = 255;
  ram[4695]  = 255;
  ram[4696]  = 255;
  ram[4697]  = 255;
  ram[4698]  = 255;
  ram[4699]  = 255;
  ram[4700]  = 255;
  ram[4701]  = 255;
  ram[4702]  = 255;
  ram[4703]  = 255;
  ram[4704]  = 255;
  ram[4705]  = 255;
  ram[4706]  = 255;
  ram[4707]  = 255;
  ram[4708]  = 255;
  ram[4709]  = 255;
  ram[4710]  = 255;
  ram[4711]  = 255;
  ram[4712]  = 255;
  ram[4713]  = 255;
  ram[4714]  = 255;
  ram[4715]  = 255;
  ram[4716]  = 255;
  ram[4717]  = 255;
  ram[4718]  = 255;
  ram[4719]  = 255;
  ram[4720]  = 255;
  ram[4721]  = 255;
  ram[4722]  = 255;
  ram[4723]  = 255;
  ram[4724]  = 255;
  ram[4725]  = 255;
  ram[4726]  = 255;
  ram[4727]  = 255;
  ram[4728]  = 255;
  ram[4729]  = 255;
  ram[4730]  = 255;
  ram[4731]  = 255;
  ram[4732]  = 255;
  ram[4733]  = 255;
  ram[4734]  = 255;
  ram[4735]  = 255;
  ram[4736]  = 255;
  ram[4737]  = 255;
  ram[4738]  = 255;
  ram[4739]  = 255;
  ram[4740]  = 255;
  ram[4741]  = 255;
  ram[4742]  = 255;
  ram[4743]  = 255;
  ram[4744]  = 255;
  ram[4745]  = 255;
  ram[4746]  = 255;
  ram[4747]  = 255;
  ram[4748]  = 255;
  ram[4749]  = 255;
  ram[4750]  = 255;
  ram[4751]  = 255;
  ram[4752]  = 255;
  ram[4753]  = 255;
  ram[4754]  = 255;
  ram[4755]  = 255;
  ram[4756]  = 255;
  ram[4757]  = 255;
  ram[4758]  = 255;
  ram[4759]  = 255;
  ram[4760]  = 255;
  ram[4761]  = 255;
  ram[4762]  = 255;
  ram[4763]  = 255;
  ram[4764]  = 255;
  ram[4765]  = 255;
  ram[4766]  = 255;
  ram[4767]  = 255;
  ram[4768]  = 255;
  ram[4769]  = 255;
  ram[4770]  = 255;
  ram[4771]  = 255;
  ram[4772]  = 255;
  ram[4773]  = 255;
  ram[4774]  = 255;
  ram[4775]  = 255;
  ram[4776]  = 255;
  ram[4777]  = 255;
  ram[4778]  = 255;
  ram[4779]  = 255;
  ram[4780]  = 255;
  ram[4781]  = 255;
  ram[4782]  = 255;
  ram[4783]  = 255;
  ram[4784]  = 255;
  ram[4785]  = 255;
  ram[4786]  = 255;
  ram[4787]  = 255;
  ram[4788]  = 255;
  ram[4789]  = 255;
  ram[4790]  = 255;
  ram[4791]  = 255;
  ram[4792]  = 255;
  ram[4793]  = 255;
  ram[4794]  = 255;
  ram[4795]  = 255;
  ram[4796]  = 255;
  ram[4797]  = 255;
  ram[4798]  = 255;
  ram[4799]  = 255;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
