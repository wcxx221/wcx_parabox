module rom_dist_g(clock, address, q);       // ROM-stored RGB bitmap for level destination
input clock;
output [7:0] q;
input [8:0] address;
reg [7:0] dout;
reg [7:0] ram [511:0];
assign q = dout;

initial begin
  ram[0]  = 255;
  ram[1]  = 255;
  ram[2]  = 255;
  ram[3]  = 255;
  ram[4]  = 255;
  ram[5]  = 255;
  ram[6]  = 255;
  ram[7]  = 162;
  ram[8]  = 162;
  ram[9]  = 162;
  ram[10]  = 162;
  ram[11]  = 162;
  ram[12]  = 255;
  ram[13]  = 255;
  ram[14]  = 255;
  ram[15]  = 255;
  ram[16]  = 255;
  ram[17]  = 255;
  ram[18]  = 255;
  ram[19]  = 255;
  ram[20]  = 255;
  ram[21]  = 255;
  ram[22]  = 255;
  ram[23]  = 255;
  ram[24]  = 255;
  ram[25]  = 162;
  ram[26]  = 162;
  ram[27]  = 162;
  ram[28]  = 162;
  ram[29]  = 162;
  ram[30]  = 162;
  ram[31]  = 162;
  ram[32]  = 162;
  ram[33]  = 162;
  ram[34]  = 255;
  ram[35]  = 255;
  ram[36]  = 255;
  ram[37]  = 255;
  ram[38]  = 255;
  ram[39]  = 255;
  ram[40]  = 255;
  ram[41]  = 255;
  ram[42]  = 255;
  ram[43]  = 162;
  ram[44]  = 162;
  ram[45]  = 162;
  ram[46]  = 162;
  ram[47]  = 162;
  ram[48]  = 162;
  ram[49]  = 162;
  ram[50]  = 162;
  ram[51]  = 162;
  ram[52]  = 162;
  ram[53]  = 162;
  ram[54]  = 162;
  ram[55]  = 162;
  ram[56]  = 255;
  ram[57]  = 255;
  ram[58]  = 255;
  ram[59]  = 255;
  ram[60]  = 255;
  ram[61]  = 255;
  ram[62]  = 162;
  ram[63]  = 162;
  ram[64]  = 162;
  ram[65]  = 162;
  ram[66]  = 162;
  ram[67]  = 162;
  ram[68]  = 162;
  ram[69]  = 162;
  ram[70]  = 162;
  ram[71]  = 162;
  ram[72]  = 162;
  ram[73]  = 162;
  ram[74]  = 162;
  ram[75]  = 162;
  ram[76]  = 162;
  ram[77]  = 255;
  ram[78]  = 255;
  ram[79]  = 255;
  ram[80]  = 255;
  ram[81]  = 255;
  ram[82]  = 162;
  ram[83]  = 162;
  ram[84]  = 162;
  ram[85]  = 162;
  ram[86]  = 162;
  ram[87]  = 162;
  ram[88]  = 162;
  ram[89]  = 162;
  ram[90]  = 162;
  ram[91]  = 162;
  ram[92]  = 162;
  ram[93]  = 162;
  ram[94]  = 162;
  ram[95]  = 162;
  ram[96]  = 162;
  ram[97]  = 255;
  ram[98]  = 255;
  ram[99]  = 255;
  ram[100]  = 255;
  ram[101]  = 162;
  ram[102]  = 162;
  ram[103]  = 162;
  ram[104]  = 162;
  ram[105]  = 162;
  ram[106]  = 162;
  ram[107]  = 162;
  ram[108]  = 255;
  ram[109]  = 255;
  ram[110]  = 255;
  ram[111]  = 162;
  ram[112]  = 162;
  ram[113]  = 162;
  ram[114]  = 162;
  ram[115]  = 162;
  ram[116]  = 162;
  ram[117]  = 162;
  ram[118]  = 255;
  ram[119]  = 255;
  ram[120]  = 255;
  ram[121]  = 162;
  ram[122]  = 162;
  ram[123]  = 162;
  ram[124]  = 162;
  ram[125]  = 162;
  ram[126]  = 255;
  ram[127]  = 255;
  ram[128]  = 255;
  ram[129]  = 255;
  ram[130]  = 255;
  ram[131]  = 255;
  ram[132]  = 255;
  ram[133]  = 162;
  ram[134]  = 162;
  ram[135]  = 162;
  ram[136]  = 162;
  ram[137]  = 162;
  ram[138]  = 255;
  ram[139]  = 255;
  ram[140]  = 162;
  ram[141]  = 162;
  ram[142]  = 162;
  ram[143]  = 162;
  ram[144]  = 162;
  ram[145]  = 162;
  ram[146]  = 255;
  ram[147]  = 255;
  ram[148]  = 255;
  ram[149]  = 255;
  ram[150]  = 255;
  ram[151]  = 255;
  ram[152]  = 255;
  ram[153]  = 162;
  ram[154]  = 162;
  ram[155]  = 162;
  ram[156]  = 162;
  ram[157]  = 162;
  ram[158]  = 162;
  ram[159]  = 255;
  ram[160]  = 162;
  ram[161]  = 162;
  ram[162]  = 162;
  ram[163]  = 162;
  ram[164]  = 162;
  ram[165]  = 255;
  ram[166]  = 255;
  ram[167]  = 255;
  ram[168]  = 255;
  ram[169]  = 255;
  ram[170]  = 255;
  ram[171]  = 255;
  ram[172]  = 255;
  ram[173]  = 255;
  ram[174]  = 162;
  ram[175]  = 162;
  ram[176]  = 162;
  ram[177]  = 162;
  ram[178]  = 162;
  ram[179]  = 255;
  ram[180]  = 162;
  ram[181]  = 162;
  ram[182]  = 162;
  ram[183]  = 162;
  ram[184]  = 162;
  ram[185]  = 255;
  ram[186]  = 255;
  ram[187]  = 255;
  ram[188]  = 255;
  ram[189]  = 255;
  ram[190]  = 255;
  ram[191]  = 255;
  ram[192]  = 255;
  ram[193]  = 255;
  ram[194]  = 162;
  ram[195]  = 162;
  ram[196]  = 162;
  ram[197]  = 162;
  ram[198]  = 162;
  ram[199]  = 255;
  ram[200]  = 162;
  ram[201]  = 162;
  ram[202]  = 162;
  ram[203]  = 162;
  ram[204]  = 162;
  ram[205]  = 255;
  ram[206]  = 255;
  ram[207]  = 255;
  ram[208]  = 255;
  ram[209]  = 255;
  ram[210]  = 255;
  ram[211]  = 255;
  ram[212]  = 255;
  ram[213]  = 255;
  ram[214]  = 162;
  ram[215]  = 162;
  ram[216]  = 162;
  ram[217]  = 162;
  ram[218]  = 162;
  ram[219]  = 255;
  ram[220]  = 162;
  ram[221]  = 162;
  ram[222]  = 162;
  ram[223]  = 162;
  ram[224]  = 162;
  ram[225]  = 255;
  ram[226]  = 255;
  ram[227]  = 255;
  ram[228]  = 255;
  ram[229]  = 255;
  ram[230]  = 255;
  ram[231]  = 255;
  ram[232]  = 255;
  ram[233]  = 255;
  ram[234]  = 162;
  ram[235]  = 162;
  ram[236]  = 162;
  ram[237]  = 162;
  ram[238]  = 162;
  ram[239]  = 255;
  ram[240]  = 162;
  ram[241]  = 162;
  ram[242]  = 162;
  ram[243]  = 162;
  ram[244]  = 162;
  ram[245]  = 162;
  ram[246]  = 255;
  ram[247]  = 255;
  ram[248]  = 255;
  ram[249]  = 255;
  ram[250]  = 255;
  ram[251]  = 255;
  ram[252]  = 255;
  ram[253]  = 162;
  ram[254]  = 162;
  ram[255]  = 162;
  ram[256]  = 162;
  ram[257]  = 162;
  ram[258]  = 162;
  ram[259]  = 255;
  ram[260]  = 255;
  ram[261]  = 162;
  ram[262]  = 162;
  ram[263]  = 162;
  ram[264]  = 162;
  ram[265]  = 162;
  ram[266]  = 255;
  ram[267]  = 255;
  ram[268]  = 255;
  ram[269]  = 255;
  ram[270]  = 255;
  ram[271]  = 255;
  ram[272]  = 255;
  ram[273]  = 162;
  ram[274]  = 162;
  ram[275]  = 162;
  ram[276]  = 162;
  ram[277]  = 162;
  ram[278]  = 255;
  ram[279]  = 255;
  ram[280]  = 255;
  ram[281]  = 162;
  ram[282]  = 162;
  ram[283]  = 162;
  ram[284]  = 162;
  ram[285]  = 162;
  ram[286]  = 162;
  ram[287]  = 162;
  ram[288]  = 255;
  ram[289]  = 255;
  ram[290]  = 255;
  ram[291]  = 162;
  ram[292]  = 162;
  ram[293]  = 162;
  ram[294]  = 162;
  ram[295]  = 162;
  ram[296]  = 162;
  ram[297]  = 162;
  ram[298]  = 255;
  ram[299]  = 255;
  ram[300]  = 255;
  ram[301]  = 255;
  ram[302]  = 162;
  ram[303]  = 162;
  ram[304]  = 162;
  ram[305]  = 162;
  ram[306]  = 162;
  ram[307]  = 162;
  ram[308]  = 162;
  ram[309]  = 162;
  ram[310]  = 162;
  ram[311]  = 162;
  ram[312]  = 162;
  ram[313]  = 162;
  ram[314]  = 162;
  ram[315]  = 162;
  ram[316]  = 162;
  ram[317]  = 255;
  ram[318]  = 255;
  ram[319]  = 255;
  ram[320]  = 255;
  ram[321]  = 255;
  ram[322]  = 162;
  ram[323]  = 162;
  ram[324]  = 162;
  ram[325]  = 162;
  ram[326]  = 162;
  ram[327]  = 162;
  ram[328]  = 162;
  ram[329]  = 162;
  ram[330]  = 162;
  ram[331]  = 162;
  ram[332]  = 162;
  ram[333]  = 162;
  ram[334]  = 162;
  ram[335]  = 162;
  ram[336]  = 162;
  ram[337]  = 255;
  ram[338]  = 255;
  ram[339]  = 255;
  ram[340]  = 255;
  ram[341]  = 255;
  ram[342]  = 255;
  ram[343]  = 162;
  ram[344]  = 162;
  ram[345]  = 162;
  ram[346]  = 162;
  ram[347]  = 162;
  ram[348]  = 162;
  ram[349]  = 162;
  ram[350]  = 162;
  ram[351]  = 162;
  ram[352]  = 162;
  ram[353]  = 162;
  ram[354]  = 162;
  ram[355]  = 162;
  ram[356]  = 255;
  ram[357]  = 255;
  ram[358]  = 255;
  ram[359]  = 255;
  ram[360]  = 255;
  ram[361]  = 255;
  ram[362]  = 255;
  ram[363]  = 255;
  ram[364]  = 255;
  ram[365]  = 162;
  ram[366]  = 162;
  ram[367]  = 162;
  ram[368]  = 162;
  ram[369]  = 162;
  ram[370]  = 162;
  ram[371]  = 162;
  ram[372]  = 162;
  ram[373]  = 162;
  ram[374]  = 255;
  ram[375]  = 255;
  ram[376]  = 255;
  ram[377]  = 255;
  ram[378]  = 255;
  ram[379]  = 255;
  ram[380]  = 255;
  ram[381]  = 255;
  ram[382]  = 255;
  ram[383]  = 255;
  ram[384]  = 255;
  ram[385]  = 255;
  ram[386]  = 255;
  ram[387]  = 162;
  ram[388]  = 162;
  ram[389]  = 162;
  ram[390]  = 162;
  ram[391]  = 162;
  ram[392]  = 255;
  ram[393]  = 255;
  ram[394]  = 255;
  ram[395]  = 255;
  ram[396]  = 255;
  ram[397]  = 255;
  ram[398]  = 255;
  ram[399]  = 255;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
