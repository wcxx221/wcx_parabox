module rom_man_r(clock, address, q);        // ROM-stored RGB bitmap for player(man)
input clock;
output [7:0] q;
input [8:0] address;
reg [7:0] dout;
reg [7:0] ram [511:0];
assign q = dout;

initial begin
  ram[0]  = 28;
  ram[1]  = 31;
  ram[2]  = 32;
  ram[3]  = 28;
  ram[4]  = 19;
  ram[5]  = 18;
  ram[6]  = 16;
  ram[7]  = 17;
  ram[8]  = 36;
  ram[9]  = 56;
  ram[10]  = 44;
  ram[11]  = 22;
  ram[12]  = 16;
  ram[13]  = 14;
  ram[14]  = 19;
  ram[15]  = 30;
  ram[16]  = 32;
  ram[17]  = 28;
  ram[18]  = 19;
  ram[19]  = 177;
  ram[20]  = 28;
  ram[21]  = 28;
  ram[22]  = 28;
  ram[23]  = 18;
  ram[24]  = 46;
  ram[25]  = 102;
  ram[26]  = 127;
  ram[27]  = 157;
  ram[28]  = 204;
  ram[29]  = 243;
  ram[30]  = 220;
  ram[31]  = 171;
  ram[32]  = 141;
  ram[33]  = 106;
  ram[34]  = 59;
  ram[35]  = 17;
  ram[36]  = 21;
  ram[37]  = 26;
  ram[38]  = 21;
  ram[39]  = 152;
  ram[40]  = 28;
  ram[41]  = 26;
  ram[42]  = 17;
  ram[43]  = 49;
  ram[44]  = 184;
  ram[45]  = 255;
  ram[46]  = 255;
  ram[47]  = 255;
  ram[48]  = 255;
  ram[49]  = 255;
  ram[50]  = 255;
  ram[51]  = 255;
  ram[52]  = 255;
  ram[53]  = 255;
  ram[54]  = 222;
  ram[55]  = 93;
  ram[56]  = 23;
  ram[57]  = 23;
  ram[58]  = 20;
  ram[59]  = 150;
  ram[60]  = 27;
  ram[61]  = 20;
  ram[62]  = 66;
  ram[63]  = 210;
  ram[64]  = 255;
  ram[65]  = 254;
  ram[66]  = 254;
  ram[67]  = 254;
  ram[68]  = 254;
  ram[69]  = 252;
  ram[70]  = 253;
  ram[71]  = 253;
  ram[72]  = 252;
  ram[73]  = 255;
  ram[74]  = 255;
  ram[75]  = 244;
  ram[76]  = 123;
  ram[77]  = 22;
  ram[78]  = 17;
  ram[79]  = 151;
  ram[80]  = 23;
  ram[81]  = 41;
  ram[82]  = 179;
  ram[83]  = 255;
  ram[84]  = 253;
  ram[85]  = 253;
  ram[86]  = 254;
  ram[87]  = 253;
  ram[88]  = 254;
  ram[89]  = 253;
  ram[90]  = 253;
  ram[91]  = 253;
  ram[92]  = 253;
  ram[93]  = 251;
  ram[94]  = 253;
  ram[95]  = 255;
  ram[96]  = 234;
  ram[97]  = 78;
  ram[98]  = 11;
  ram[99]  = 151;
  ram[100]  = 17;
  ram[101]  = 93;
  ram[102]  = 239;
  ram[103]  = 255;
  ram[104]  = 252;
  ram[105]  = 254;
  ram[106]  = 251;
  ram[107]  = 251;
  ram[108]  = 252;
  ram[109]  = 251;
  ram[110]  = 253;
  ram[111]  = 255;
  ram[112]  = 255;
  ram[113]  = 250;
  ram[114]  = 251;
  ram[115]  = 255;
  ram[116]  = 255;
  ram[117]  = 165;
  ram[118]  = 24;
  ram[119]  = 148;
  ram[120]  = 18;
  ram[121]  = 136;
  ram[122]  = 255;
  ram[123]  = 255;
  ram[124]  = 253;
  ram[125]  = 251;
  ram[126]  = 254;
  ram[127]  = 255;
  ram[128]  = 254;
  ram[129]  = 250;
  ram[130]  = 251;
  ram[131]  = 255;
  ram[132]  = 255;
  ram[133]  = 250;
  ram[134]  = 251;
  ram[135]  = 255;
  ram[136]  = 255;
  ram[137]  = 213;
  ram[138]  = 47;
  ram[139]  = 144;
  ram[140]  = 22;
  ram[141]  = 156;
  ram[142]  = 253;
  ram[143]  = 243;
  ram[144]  = 233;
  ram[145]  = 226;
  ram[146]  = 215;
  ram[147]  = 209;
  ram[148]  = 223;
  ram[149]  = 226;
  ram[150]  = 219;
  ram[151]  = 203;
  ram[152]  = 204;
  ram[153]  = 218;
  ram[154]  = 226;
  ram[155]  = 234;
  ram[156]  = 244;
  ram[157]  = 226;
  ram[158]  = 56;
  ram[159]  = 143;
  ram[160]  = 24;
  ram[161]  = 137;
  ram[162]  = 227;
  ram[163]  = 216;
  ram[164]  = 229;
  ram[165]  = 210;
  ram[166]  = 94;
  ram[167]  = 68;
  ram[168]  = 179;
  ram[169]  = 252;
  ram[170]  = 205;
  ram[171]  = 71;
  ram[172]  = 69;
  ram[173]  = 184;
  ram[174]  = 241;
  ram[175]  = 221;
  ram[176]  = 216;
  ram[177]  = 215;
  ram[178]  = 61;
  ram[179]  = 143;
  ram[180]  = 21;
  ram[181]  = 98;
  ram[182]  = 203;
  ram[183]  = 244;
  ram[184]  = 255;
  ram[185]  = 191;
  ram[186]  = 51;
  ram[187]  = 43;
  ram[188]  = 150;
  ram[189]  = 255;
  ram[190]  = 193;
  ram[191]  = 45;
  ram[192]  = 36;
  ram[193]  = 159;
  ram[194]  = 255;
  ram[195]  = 255;
  ram[196]  = 230;
  ram[197]  = 185;
  ram[198]  = 53;
  ram[199]  = 146;
  ram[200]  = 27;
  ram[201]  = 29;
  ram[202]  = 68;
  ram[203]  = 153;
  ram[204]  = 251;
  ram[205]  = 229;
  ram[206]  = 75;
  ram[207]  = 57;
  ram[208]  = 195;
  ram[209]  = 255;
  ram[210]  = 222;
  ram[211]  = 76;
  ram[212]  = 52;
  ram[213]  = 197;
  ram[214]  = 255;
  ram[215]  = 211;
  ram[216]  = 105;
  ram[217]  = 54;
  ram[218]  = 21;
  ram[219]  = 151;
  ram[220]  = 31;
  ram[221]  = 25;
  ram[222]  = 16;
  ram[223]  = 15;
  ram[224]  = 117;
  ram[225]  = 249;
  ram[226]  = 205;
  ram[227]  = 185;
  ram[228]  = 249;
  ram[229]  = 255;
  ram[230]  = 254;
  ram[231]  = 202;
  ram[232]  = 189;
  ram[233]  = 255;
  ram[234]  = 198;
  ram[235]  = 60;
  ram[236]  = 7;
  ram[237]  = 20;
  ram[238]  = 21;
  ram[239]  = 151;
  ram[240]  = 28;
  ram[241]  = 26;
  ram[242]  = 24;
  ram[243]  = 24;
  ram[244]  = 33;
  ram[245]  = 172;
  ram[246]  = 255;
  ram[247]  = 255;
  ram[248]  = 254;
  ram[249]  = 253;
  ram[250]  = 252;
  ram[251]  = 255;
  ram[252]  = 255;
  ram[253]  = 218;
  ram[254]  = 69;
  ram[255]  = 18;
  ram[256]  = 28;
  ram[257]  = 24;
  ram[258]  = 21;
  ram[259]  = 151;
  ram[260]  = 28;
  ram[261]  = 25;
  ram[262]  = 30;
  ram[263]  = 29;
  ram[264]  = 20;
  ram[265]  = 47;
  ram[266]  = 144;
  ram[267]  = 222;
  ram[268]  = 250;
  ram[269]  = 254;
  ram[270]  = 249;
  ram[271]  = 240;
  ram[272]  = 183;
  ram[273]  = 75;
  ram[274]  = 21;
  ram[275]  = 25;
  ram[276]  = 32;
  ram[277]  = 23;
  ram[278]  = 19;
  ram[279]  = 151;
  ram[280]  = 31;
  ram[281]  = 26;
  ram[282]  = 27;
  ram[283]  = 29;
  ram[284]  = 29;
  ram[285]  = 22;
  ram[286]  = 26;
  ram[287]  = 55;
  ram[288]  = 98;
  ram[289]  = 115;
  ram[290]  = 105;
  ram[291]  = 77;
  ram[292]  = 38;
  ram[293]  = 24;
  ram[294]  = 22;
  ram[295]  = 27;
  ram[296]  = 28;
  ram[297]  = 25;
  ram[298]  = 20;
  ram[299]  = 151;
  ram[300]  = 29;
  ram[301]  = 18;
  ram[302]  = 61;
  ram[303]  = 182;
  ram[304]  = 184;
  ram[305]  = 64;
  ram[306]  = 28;
  ram[307]  = 27;
  ram[308]  = 24;
  ram[309]  = 28;
  ram[310]  = 26;
  ram[311]  = 25;
  ram[312]  = 30;
  ram[313]  = 32;
  ram[314]  = 105;
  ram[315]  = 194;
  ram[316]  = 134;
  ram[317]  = 29;
  ram[318]  = 18;
  ram[319]  = 151;
  ram[320]  = 28;
  ram[321]  = 16;
  ram[322]  = 80;
  ram[323]  = 246;
  ram[324]  = 244;
  ram[325]  = 83;
  ram[326]  = 23;
  ram[327]  = 33;
  ram[328]  = 33;
  ram[329]  = 32;
  ram[330]  = 33;
  ram[331]  = 35;
  ram[332]  = 36;
  ram[333]  = 37;
  ram[334]  = 157;
  ram[335]  = 255;
  ram[336]  = 175;
  ram[337]  = 33;
  ram[338]  = 16;
  ram[339]  = 151;
  ram[340]  = 28;
  ram[341]  = 25;
  ram[342]  = 30;
  ram[343]  = 66;
  ram[344]  = 63;
  ram[345]  = 31;
  ram[346]  = 50;
  ram[347]  = 60;
  ram[348]  = 54;
  ram[349]  = 41;
  ram[350]  = 45;
  ram[351]  = 56;
  ram[352]  = 57;
  ram[353]  = 43;
  ram[354]  = 38;
  ram[355]  = 71;
  ram[356]  = 49;
  ram[357]  = 25;
  ram[358]  = 20;
  ram[359]  = 151;
  ram[360]  = 30;
  ram[361]  = 27;
  ram[362]  = 25;
  ram[363]  = 20;
  ram[364]  = 19;
  ram[365]  = 43;
  ram[366]  = 71;
  ram[367]  = 76;
  ram[368]  = 71;
  ram[369]  = 48;
  ram[370]  = 55;
  ram[371]  = 71;
  ram[372]  = 71;
  ram[373]  = 62;
  ram[374]  = 30;
  ram[375]  = 13;
  ram[376]  = 27;
  ram[377]  = 28;
  ram[378]  = 20;
  ram[379]  = 151;
  ram[380]  = 28;
  ram[381]  = 29;
  ram[382]  = 29;
  ram[383]  = 29;
  ram[384]  = 28;
  ram[385]  = 33;
  ram[386]  = 41;
  ram[387]  = 39;
  ram[388]  = 39;
  ram[389]  = 32;
  ram[390]  = 38;
  ram[391]  = 42;
  ram[392]  = 38;
  ram[393]  = 36;
  ram[394]  = 29;
  ram[395]  = 28;
  ram[396]  = 28;
  ram[397]  = 27;
  ram[398]  = 21;
  ram[399]  = 151;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
