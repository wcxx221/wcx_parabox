module rom_cai_g(clock, address, q);        // ROM-stored RGB bitmap for cai
input clock;
output [7:0] q;
input [8:0] address;
reg [7:0] dout;
reg [7:0] ram [511:0];
assign q = dout;

initial begin
  ram[0]  = 255;
  ram[1]  = 255;
  ram[2]  = 255;
  ram[3]  = 255;
  ram[4]  = 255;
  ram[5]  = 255;
  ram[6]  = 255;
  ram[7]  = 255;
  ram[8]  = 255;
  ram[9]  = 72;
  ram[10]  = 72;
  ram[11]  = 255;
  ram[12]  = 255;
  ram[13]  = 255;
  ram[14]  = 255;
  ram[15]  = 255;
  ram[16]  = 255;
  ram[17]  = 255;
  ram[18]  = 255;
  ram[19]  = 255;
  ram[20]  = 255;
  ram[21]  = 255;
  ram[22]  = 255;
  ram[23]  = 255;
  ram[24]  = 255;
  ram[25]  = 255;
  ram[26]  = 255;
  ram[27]  = 255;
  ram[28]  = 72;
  ram[29]  = 72;
  ram[30]  = 72;
  ram[31]  = 72;
  ram[32]  = 255;
  ram[33]  = 255;
  ram[34]  = 255;
  ram[35]  = 255;
  ram[36]  = 255;
  ram[37]  = 255;
  ram[38]  = 255;
  ram[39]  = 255;
  ram[40]  = 255;
  ram[41]  = 255;
  ram[42]  = 255;
  ram[43]  = 255;
  ram[44]  = 255;
  ram[45]  = 255;
  ram[46]  = 255;
  ram[47]  = 72;
  ram[48]  = 72;
  ram[49]  = 72;
  ram[50]  = 72;
  ram[51]  = 72;
  ram[52]  = 72;
  ram[53]  = 255;
  ram[54]  = 255;
  ram[55]  = 255;
  ram[56]  = 255;
  ram[57]  = 255;
  ram[58]  = 255;
  ram[59]  = 255;
  ram[60]  = 255;
  ram[61]  = 255;
  ram[62]  = 255;
  ram[63]  = 255;
  ram[64]  = 255;
  ram[65]  = 255;
  ram[66]  = 255;
  ram[67]  = 72;
  ram[68]  = 72;
  ram[69]  = 72;
  ram[70]  = 72;
  ram[71]  = 72;
  ram[72]  = 72;
  ram[73]  = 255;
  ram[74]  = 255;
  ram[75]  = 255;
  ram[76]  = 255;
  ram[77]  = 255;
  ram[78]  = 255;
  ram[79]  = 255;
  ram[80]  = 255;
  ram[81]  = 255;
  ram[82]  = 255;
  ram[83]  = 255;
  ram[84]  = 255;
  ram[85]  = 255;
  ram[86]  = 72;
  ram[87]  = 72;
  ram[88]  = 72;
  ram[89]  = 72;
  ram[90]  = 72;
  ram[91]  = 72;
  ram[92]  = 72;
  ram[93]  = 72;
  ram[94]  = 255;
  ram[95]  = 255;
  ram[96]  = 255;
  ram[97]  = 255;
  ram[98]  = 255;
  ram[99]  = 255;
  ram[100]  = 255;
  ram[101]  = 255;
  ram[102]  = 255;
  ram[103]  = 255;
  ram[104]  = 255;
  ram[105]  = 255;
  ram[106]  = 72;
  ram[107]  = 72;
  ram[108]  = 72;
  ram[109]  = 72;
  ram[110]  = 72;
  ram[111]  = 72;
  ram[112]  = 72;
  ram[113]  = 72;
  ram[114]  = 255;
  ram[115]  = 255;
  ram[116]  = 255;
  ram[117]  = 255;
  ram[118]  = 255;
  ram[119]  = 255;
  ram[120]  = 255;
  ram[121]  = 255;
  ram[122]  = 255;
  ram[123]  = 255;
  ram[124]  = 255;
  ram[125]  = 72;
  ram[126]  = 72;
  ram[127]  = 72;
  ram[128]  = 72;
  ram[129]  = 72;
  ram[130]  = 72;
  ram[131]  = 72;
  ram[132]  = 72;
  ram[133]  = 72;
  ram[134]  = 72;
  ram[135]  = 255;
  ram[136]  = 255;
  ram[137]  = 255;
  ram[138]  = 255;
  ram[139]  = 255;
  ram[140]  = 255;
  ram[141]  = 255;
  ram[142]  = 255;
  ram[143]  = 255;
  ram[144]  = 255;
  ram[145]  = 72;
  ram[146]  = 72;
  ram[147]  = 72;
  ram[148]  = 72;
  ram[149]  = 72;
  ram[150]  = 72;
  ram[151]  = 72;
  ram[152]  = 72;
  ram[153]  = 72;
  ram[154]  = 72;
  ram[155]  = 255;
  ram[156]  = 255;
  ram[157]  = 255;
  ram[158]  = 255;
  ram[159]  = 255;
  ram[160]  = 255;
  ram[161]  = 255;
  ram[162]  = 255;
  ram[163]  = 255;
  ram[164]  = 72;
  ram[165]  = 72;
  ram[166]  = 72;
  ram[167]  = 72;
  ram[168]  = 72;
  ram[169]  = 72;
  ram[170]  = 72;
  ram[171]  = 72;
  ram[172]  = 72;
  ram[173]  = 72;
  ram[174]  = 72;
  ram[175]  = 72;
  ram[176]  = 255;
  ram[177]  = 255;
  ram[178]  = 255;
  ram[179]  = 255;
  ram[180]  = 255;
  ram[181]  = 255;
  ram[182]  = 255;
  ram[183]  = 255;
  ram[184]  = 72;
  ram[185]  = 72;
  ram[186]  = 72;
  ram[187]  = 72;
  ram[188]  = 72;
  ram[189]  = 255;
  ram[190]  = 255;
  ram[191]  = 72;
  ram[192]  = 72;
  ram[193]  = 72;
  ram[194]  = 72;
  ram[195]  = 72;
  ram[196]  = 255;
  ram[197]  = 255;
  ram[198]  = 255;
  ram[199]  = 255;
  ram[200]  = 255;
  ram[201]  = 255;
  ram[202]  = 255;
  ram[203]  = 72;
  ram[204]  = 72;
  ram[205]  = 72;
  ram[206]  = 72;
  ram[207]  = 72;
  ram[208]  = 72;
  ram[209]  = 255;
  ram[210]  = 255;
  ram[211]  = 72;
  ram[212]  = 72;
  ram[213]  = 72;
  ram[214]  = 72;
  ram[215]  = 72;
  ram[216]  = 72;
  ram[217]  = 255;
  ram[218]  = 255;
  ram[219]  = 255;
  ram[220]  = 255;
  ram[221]  = 255;
  ram[222]  = 255;
  ram[223]  = 72;
  ram[224]  = 72;
  ram[225]  = 72;
  ram[226]  = 72;
  ram[227]  = 72;
  ram[228]  = 255;
  ram[229]  = 255;
  ram[230]  = 255;
  ram[231]  = 255;
  ram[232]  = 72;
  ram[233]  = 72;
  ram[234]  = 72;
  ram[235]  = 72;
  ram[236]  = 72;
  ram[237]  = 255;
  ram[238]  = 255;
  ram[239]  = 255;
  ram[240]  = 255;
  ram[241]  = 255;
  ram[242]  = 72;
  ram[243]  = 72;
  ram[244]  = 72;
  ram[245]  = 72;
  ram[246]  = 72;
  ram[247]  = 72;
  ram[248]  = 255;
  ram[249]  = 255;
  ram[250]  = 255;
  ram[251]  = 255;
  ram[252]  = 72;
  ram[253]  = 72;
  ram[254]  = 72;
  ram[255]  = 72;
  ram[256]  = 72;
  ram[257]  = 72;
  ram[258]  = 255;
  ram[259]  = 255;
  ram[260]  = 255;
  ram[261]  = 255;
  ram[262]  = 72;
  ram[263]  = 72;
  ram[264]  = 72;
  ram[265]  = 72;
  ram[266]  = 72;
  ram[267]  = 255;
  ram[268]  = 255;
  ram[269]  = 255;
  ram[270]  = 255;
  ram[271]  = 255;
  ram[272]  = 255;
  ram[273]  = 72;
  ram[274]  = 72;
  ram[275]  = 72;
  ram[276]  = 72;
  ram[277]  = 72;
  ram[278]  = 255;
  ram[279]  = 255;
  ram[280]  = 255;
  ram[281]  = 72;
  ram[282]  = 72;
  ram[283]  = 72;
  ram[284]  = 72;
  ram[285]  = 72;
  ram[286]  = 72;
  ram[287]  = 255;
  ram[288]  = 255;
  ram[289]  = 255;
  ram[290]  = 255;
  ram[291]  = 255;
  ram[292]  = 255;
  ram[293]  = 72;
  ram[294]  = 72;
  ram[295]  = 72;
  ram[296]  = 72;
  ram[297]  = 72;
  ram[298]  = 72;
  ram[299]  = 255;
  ram[300]  = 255;
  ram[301]  = 72;
  ram[302]  = 72;
  ram[303]  = 72;
  ram[304]  = 72;
  ram[305]  = 72;
  ram[306]  = 72;
  ram[307]  = 72;
  ram[308]  = 72;
  ram[309]  = 72;
  ram[310]  = 72;
  ram[311]  = 72;
  ram[312]  = 72;
  ram[313]  = 72;
  ram[314]  = 72;
  ram[315]  = 72;
  ram[316]  = 72;
  ram[317]  = 72;
  ram[318]  = 72;
  ram[319]  = 255;
  ram[320]  = 72;
  ram[321]  = 72;
  ram[322]  = 72;
  ram[323]  = 72;
  ram[324]  = 72;
  ram[325]  = 72;
  ram[326]  = 72;
  ram[327]  = 72;
  ram[328]  = 72;
  ram[329]  = 72;
  ram[330]  = 72;
  ram[331]  = 72;
  ram[332]  = 72;
  ram[333]  = 72;
  ram[334]  = 72;
  ram[335]  = 72;
  ram[336]  = 72;
  ram[337]  = 72;
  ram[338]  = 72;
  ram[339]  = 72;
  ram[340]  = 72;
  ram[341]  = 72;
  ram[342]  = 72;
  ram[343]  = 72;
  ram[344]  = 72;
  ram[345]  = 72;
  ram[346]  = 72;
  ram[347]  = 72;
  ram[348]  = 72;
  ram[349]  = 72;
  ram[350]  = 72;
  ram[351]  = 72;
  ram[352]  = 72;
  ram[353]  = 72;
  ram[354]  = 72;
  ram[355]  = 72;
  ram[356]  = 72;
  ram[357]  = 72;
  ram[358]  = 72;
  ram[359]  = 72;
  ram[360]  = 72;
  ram[361]  = 72;
  ram[362]  = 72;
  ram[363]  = 72;
  ram[364]  = 72;
  ram[365]  = 72;
  ram[366]  = 72;
  ram[367]  = 72;
  ram[368]  = 72;
  ram[369]  = 72;
  ram[370]  = 72;
  ram[371]  = 72;
  ram[372]  = 72;
  ram[373]  = 72;
  ram[374]  = 72;
  ram[375]  = 72;
  ram[376]  = 72;
  ram[377]  = 72;
  ram[378]  = 72;
  ram[379]  = 72;
  ram[380]  = 255;
  ram[381]  = 72;
  ram[382]  = 72;
  ram[383]  = 72;
  ram[384]  = 72;
  ram[385]  = 72;
  ram[386]  = 72;
  ram[387]  = 72;
  ram[388]  = 72;
  ram[389]  = 72;
  ram[390]  = 72;
  ram[391]  = 72;
  ram[392]  = 72;
  ram[393]  = 72;
  ram[394]  = 72;
  ram[395]  = 72;
  ram[396]  = 72;
  ram[397]  = 72;
  ram[398]  = 72;
  ram[399]  = 255;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
