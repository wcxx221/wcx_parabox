module rom_cai(clock, address, q);     // ROM-stored RGB bitmap for cai_dan
input clock;
output [7:0] q;
input [11:0] address;
reg [7:0] dout;
reg [7:0] ram [4095:0];
assign q = dout;

initial begin
  ram[0]  = 255;
  ram[1]  = 255;
  ram[2]  = 255;
  ram[3]  = 255;
  ram[4]  = 255;
  ram[5]  = 255;
  ram[6]  = 255;
  ram[7]  = 255;
  ram[8]  = 255;
  ram[9]  = 255;
  ram[10]  = 255;
  ram[11]  = 255;
  ram[12]  = 255;
  ram[13]  = 255;
  ram[14]  = 255;
  ram[15]  = 255;
  ram[16]  = 255;
  ram[17]  = 255;
  ram[18]  = 255;
  ram[19]  = 255;
  ram[20]  = 255;
  ram[21]  = 255;
  ram[22]  = 255;
  ram[23]  = 255;
  ram[24]  = 255;
  ram[25]  = 255;
  ram[26]  = 255;
  ram[27]  = 255;
  ram[28]  = 255;
  ram[29]  = 255;
  ram[30]  = 255;
  ram[31]  = 255;
  ram[32]  = 255;
  ram[33]  = 255;
  ram[34]  = 255;
  ram[35]  = 255;
  ram[36]  = 255;
  ram[37]  = 255;
  ram[38]  = 255;
  ram[39]  = 255;
  ram[40]  = 255;
  ram[41]  = 255;
  ram[42]  = 255;
  ram[43]  = 255;
  ram[44]  = 255;
  ram[45]  = 255;
  ram[46]  = 255;
  ram[47]  = 255;
  ram[48]  = 255;
  ram[49]  = 255;
  ram[50]  = 255;
  ram[51]  = 255;
  ram[52]  = 255;
  ram[53]  = 255;
  ram[54]  = 255;
  ram[55]  = 255;
  ram[56]  = 255;
  ram[57]  = 255;
  ram[58]  = 255;
  ram[59]  = 255;
  ram[60]  = 255;
  ram[61]  = 255;
  ram[62]  = 255;
  ram[63]  = 255;
  ram[64]  = 255;
  ram[65]  = 255;
  ram[66]  = 255;
  ram[67]  = 255;
  ram[68]  = 255;
  ram[69]  = 255;
  ram[70]  = 255;
  ram[71]  = 255;
  ram[72]  = 255;
  ram[73]  = 255;
  ram[74]  = 255;
  ram[75]  = 255;
  ram[76]  = 255;
  ram[77]  = 255;
  ram[78]  = 255;
  ram[79]  = 255;
  ram[80]  = 255;
  ram[81]  = 255;
  ram[82]  = 255;
  ram[83]  = 255;
  ram[84]  = 255;
  ram[85]  = 255;
  ram[86]  = 255;
  ram[87]  = 255;
  ram[88]  = 255;
  ram[89]  = 255;
  ram[90]  = 255;
  ram[91]  = 255;
  ram[92]  = 255;
  ram[93]  = 255;
  ram[94]  = 255;
  ram[95]  = 255;
  ram[96]  = 255;
  ram[97]  = 255;
  ram[98]  = 255;
  ram[99]  = 255;
  ram[100]  = 255;
  ram[101]  = 255;
  ram[102]  = 255;
  ram[103]  = 255;
  ram[104]  = 255;
  ram[105]  = 255;
  ram[106]  = 255;
  ram[107]  = 255;
  ram[108]  = 255;
  ram[109]  = 255;
  ram[110]  = 255;
  ram[111]  = 255;
  ram[112]  = 255;
  ram[113]  = 255;
  ram[114]  = 255;
  ram[115]  = 255;
  ram[116]  = 255;
  ram[117]  = 255;
  ram[118]  = 255;
  ram[119]  = 255;
  ram[120]  = 255;
  ram[121]  = 255;
  ram[122]  = 255;
  ram[123]  = 255;
  ram[124]  = 255;
  ram[125]  = 255;
  ram[126]  = 255;
  ram[127]  = 255;
  ram[128]  = 255;
  ram[129]  = 255;
  ram[130]  = 255;
  ram[131]  = 255;
  ram[132]  = 255;
  ram[133]  = 255;
  ram[134]  = 255;
  ram[135]  = 255;
  ram[136]  = 255;
  ram[137]  = 255;
  ram[138]  = 255;
  ram[139]  = 255;
  ram[140]  = 255;
  ram[141]  = 255;
  ram[142]  = 255;
  ram[143]  = 255;
  ram[144]  = 255;
  ram[145]  = 255;
  ram[146]  = 255;
  ram[147]  = 255;
  ram[148]  = 255;
  ram[149]  = 255;
  ram[150]  = 255;
  ram[151]  = 255;
  ram[152]  = 255;
  ram[153]  = 255;
  ram[154]  = 255;
  ram[155]  = 255;
  ram[156]  = 255;
  ram[157]  = 255;
  ram[158]  = 255;
  ram[159]  = 255;
  ram[160]  = 255;
  ram[161]  = 255;
  ram[162]  = 255;
  ram[163]  = 255;
  ram[164]  = 255;
  ram[165]  = 255;
  ram[166]  = 255;
  ram[167]  = 255;
  ram[168]  = 255;
  ram[169]  = 255;
  ram[170]  = 255;
  ram[171]  = 255;
  ram[172]  = 255;
  ram[173]  = 255;
  ram[174]  = 255;
  ram[175]  = 255;
  ram[176]  = 255;
  ram[177]  = 255;
  ram[178]  = 255;
  ram[179]  = 255;
  ram[180]  = 255;
  ram[181]  = 255;
  ram[182]  = 255;
  ram[183]  = 255;
  ram[184]  = 255;
  ram[185]  = 255;
  ram[186]  = 255;
  ram[187]  = 255;
  ram[188]  = 255;
  ram[189]  = 255;
  ram[190]  = 255;
  ram[191]  = 255;
  ram[192]  = 255;
  ram[193]  = 255;
  ram[194]  = 255;
  ram[195]  = 255;
  ram[196]  = 255;
  ram[197]  = 255;
  ram[198]  = 255;
  ram[199]  = 255;
  ram[200]  = 255;
  ram[201]  = 255;
  ram[202]  = 255;
  ram[203]  = 255;
  ram[204]  = 255;
  ram[205]  = 255;
  ram[206]  = 255;
  ram[207]  = 255;
  ram[208]  = 255;
  ram[209]  = 255;
  ram[210]  = 255;
  ram[211]  = 255;
  ram[212]  = 255;
  ram[213]  = 255;
  ram[214]  = 255;
  ram[215]  = 255;
  ram[216]  = 255;
  ram[217]  = 255;
  ram[218]  = 255;
  ram[219]  = 255;
  ram[220]  = 255;
  ram[221]  = 255;
  ram[222]  = 255;
  ram[223]  = 255;
  ram[224]  = 255;
  ram[225]  = 255;
  ram[226]  = 255;
  ram[227]  = 255;
  ram[228]  = 255;
  ram[229]  = 255;
  ram[230]  = 255;
  ram[231]  = 255;
  ram[232]  = 255;
  ram[233]  = 255;
  ram[234]  = 255;
  ram[235]  = 255;
  ram[236]  = 255;
  ram[237]  = 255;
  ram[238]  = 255;
  ram[239]  = 255;
  ram[240]  = 255;
  ram[241]  = 255;
  ram[242]  = 255;
  ram[243]  = 255;
  ram[244]  = 255;
  ram[245]  = 255;
  ram[246]  = 255;
  ram[247]  = 255;
  ram[248]  = 255;
  ram[249]  = 255;
  ram[250]  = 255;
  ram[251]  = 255;
  ram[252]  = 255;
  ram[253]  = 255;
  ram[254]  = 255;
  ram[255]  = 255;
  ram[256]  = 255;
  ram[257]  = 255;
  ram[258]  = 255;
  ram[259]  = 255;
  ram[260]  = 255;
  ram[261]  = 255;
  ram[262]  = 255;
  ram[263]  = 255;
  ram[264]  = 255;
  ram[265]  = 255;
  ram[266]  = 255;
  ram[267]  = 255;
  ram[268]  = 255;
  ram[269]  = 255;
  ram[270]  = 255;
  ram[271]  = 255;
  ram[272]  = 255;
  ram[273]  = 255;
  ram[274]  = 255;
  ram[275]  = 255;
  ram[276]  = 255;
  ram[277]  = 255;
  ram[278]  = 255;
  ram[279]  = 255;
  ram[280]  = 255;
  ram[281]  = 255;
  ram[282]  = 255;
  ram[283]  = 255;
  ram[284]  = 255;
  ram[285]  = 255;
  ram[286]  = 255;
  ram[287]  = 255;
  ram[288]  = 255;
  ram[289]  = 255;
  ram[290]  = 255;
  ram[291]  = 255;
  ram[292]  = 255;
  ram[293]  = 255;
  ram[294]  = 255;
  ram[295]  = 255;
  ram[296]  = 255;
  ram[297]  = 255;
  ram[298]  = 255;
  ram[299]  = 255;
  ram[300]  = 255;
  ram[301]  = 255;
  ram[302]  = 255;
  ram[303]  = 255;
  ram[304]  = 255;
  ram[305]  = 255;
  ram[306]  = 255;
  ram[307]  = 255;
  ram[308]  = 255;
  ram[309]  = 255;
  ram[310]  = 255;
  ram[311]  = 255;
  ram[312]  = 255;
  ram[313]  = 255;
  ram[314]  = 255;
  ram[315]  = 255;
  ram[316]  = 255;
  ram[317]  = 255;
  ram[318]  = 255;
  ram[319]  = 255;
  ram[320]  = 255;
  ram[321]  = 255;
  ram[322]  = 255;
  ram[323]  = 255;
  ram[324]  = 255;
  ram[325]  = 255;
  ram[326]  = 255;
  ram[327]  = 255;
  ram[328]  = 255;
  ram[329]  = 255;
  ram[330]  = 255;
  ram[331]  = 255;
  ram[332]  = 255;
  ram[333]  = 255;
  ram[334]  = 255;
  ram[335]  = 255;
  ram[336]  = 255;
  ram[337]  = 255;
  ram[338]  = 255;
  ram[339]  = 255;
  ram[340]  = 255;
  ram[341]  = 255;
  ram[342]  = 255;
  ram[343]  = 255;
  ram[344]  = 255;
  ram[345]  = 255;
  ram[346]  = 255;
  ram[347]  = 255;
  ram[348]  = 255;
  ram[349]  = 255;
  ram[350]  = 255;
  ram[351]  = 255;
  ram[352]  = 255;
  ram[353]  = 255;
  ram[354]  = 255;
  ram[355]  = 255;
  ram[356]  = 255;
  ram[357]  = 255;
  ram[358]  = 255;
  ram[359]  = 255;
  ram[360]  = 255;
  ram[361]  = 255;
  ram[362]  = 255;
  ram[363]  = 255;
  ram[364]  = 255;
  ram[365]  = 255;
  ram[366]  = 255;
  ram[367]  = 255;
  ram[368]  = 255;
  ram[369]  = 255;
  ram[370]  = 255;
  ram[371]  = 255;
  ram[372]  = 255;
  ram[373]  = 255;
  ram[374]  = 255;
  ram[375]  = 255;
  ram[376]  = 255;
  ram[377]  = 255;
  ram[378]  = 255;
  ram[379]  = 255;
  ram[380]  = 255;
  ram[381]  = 255;
  ram[382]  = 255;
  ram[383]  = 255;
  ram[384]  = 255;
  ram[385]  = 255;
  ram[386]  = 255;
  ram[387]  = 255;
  ram[388]  = 255;
  ram[389]  = 255;
  ram[390]  = 255;
  ram[391]  = 255;
  ram[392]  = 255;
  ram[393]  = 255;
  ram[394]  = 255;
  ram[395]  = 255;
  ram[396]  = 255;
  ram[397]  = 255;
  ram[398]  = 255;
  ram[399]  = 255;
  ram[400]  = 255;
  ram[401]  = 255;
  ram[402]  = 255;
  ram[403]  = 255;
  ram[404]  = 255;
  ram[405]  = 255;
  ram[406]  = 255;
  ram[407]  = 255;
  ram[408]  = 255;
  ram[409]  = 255;
  ram[410]  = 255;
  ram[411]  = 255;
  ram[412]  = 255;
  ram[413]  = 255;
  ram[414]  = 255;
  ram[415]  = 255;
  ram[416]  = 255;
  ram[417]  = 255;
  ram[418]  = 255;
  ram[419]  = 255;
  ram[420]  = 255;
  ram[421]  = 255;
  ram[422]  = 255;
  ram[423]  = 255;
  ram[424]  = 255;
  ram[425]  = 255;
  ram[426]  = 255;
  ram[427]  = 255;
  ram[428]  = 255;
  ram[429]  = 255;
  ram[430]  = 255;
  ram[431]  = 255;
  ram[432]  = 255;
  ram[433]  = 255;
  ram[434]  = 255;
  ram[435]  = 255;
  ram[436]  = 255;
  ram[437]  = 255;
  ram[438]  = 255;
  ram[439]  = 255;
  ram[440]  = 255;
  ram[441]  = 255;
  ram[442]  = 255;
  ram[443]  = 255;
  ram[444]  = 255;
  ram[445]  = 255;
  ram[446]  = 255;
  ram[447]  = 255;
  ram[448]  = 255;
  ram[449]  = 255;
  ram[450]  = 255;
  ram[451]  = 255;
  ram[452]  = 255;
  ram[453]  = 255;
  ram[454]  = 255;
  ram[455]  = 255;
  ram[456]  = 255;
  ram[457]  = 255;
  ram[458]  = 255;
  ram[459]  = 255;
  ram[460]  = 255;
  ram[461]  = 255;
  ram[462]  = 255;
  ram[463]  = 255;
  ram[464]  = 255;
  ram[465]  = 255;
  ram[466]  = 255;
  ram[467]  = 255;
  ram[468]  = 255;
  ram[469]  = 255;
  ram[470]  = 255;
  ram[471]  = 255;
  ram[472]  = 255;
  ram[473]  = 255;
  ram[474]  = 255;
  ram[475]  = 255;
  ram[476]  = 255;
  ram[477]  = 255;
  ram[478]  = 255;
  ram[479]  = 255;
  ram[480]  = 255;
  ram[481]  = 255;
  ram[482]  = 255;
  ram[483]  = 255;
  ram[484]  = 255;
  ram[485]  = 255;
  ram[486]  = 255;
  ram[487]  = 255;
  ram[488]  = 255;
  ram[489]  = 255;
  ram[490]  = 255;
  ram[491]  = 255;
  ram[492]  = 255;
  ram[493]  = 255;
  ram[494]  = 255;
  ram[495]  = 255;
  ram[496]  = 255;
  ram[497]  = 255;
  ram[498]  = 255;
  ram[499]  = 255;
  ram[500]  = 255;
  ram[501]  = 255;
  ram[502]  = 255;
  ram[503]  = 255;
  ram[504]  = 255;
  ram[505]  = 255;
  ram[506]  = 255;
  ram[507]  = 255;
  ram[508]  = 255;
  ram[509]  = 255;
  ram[510]  = 255;
  ram[511]  = 255;
  ram[512]  = 255;
  ram[513]  = 255;
  ram[514]  = 255;
  ram[515]  = 255;
  ram[516]  = 255;
  ram[517]  = 255;
  ram[518]  = 255;
  ram[519]  = 255;
  ram[520]  = 255;
  ram[521]  = 255;
  ram[522]  = 255;
  ram[523]  = 255;
  ram[524]  = 255;
  ram[525]  = 255;
  ram[526]  = 255;
  ram[527]  = 255;
  ram[528]  = 255;
  ram[529]  = 255;
  ram[530]  = 255;
  ram[531]  = 255;
  ram[532]  = 255;
  ram[533]  = 255;
  ram[534]  = 255;
  ram[535]  = 255;
  ram[536]  = 255;
  ram[537]  = 255;
  ram[538]  = 255;
  ram[539]  = 255;
  ram[540]  = 255;
  ram[541]  = 255;
  ram[542]  = 255;
  ram[543]  = 255;
  ram[544]  = 255;
  ram[545]  = 255;
  ram[546]  = 255;
  ram[547]  = 255;
  ram[548]  = 255;
  ram[549]  = 255;
  ram[550]  = 255;
  ram[551]  = 255;
  ram[552]  = 255;
  ram[553]  = 255;
  ram[554]  = 255;
  ram[555]  = 255;
  ram[556]  = 255;
  ram[557]  = 255;
  ram[558]  = 255;
  ram[559]  = 255;
  ram[560]  = 255;
  ram[561]  = 255;
  ram[562]  = 255;
  ram[563]  = 255;
  ram[564]  = 255;
  ram[565]  = 255;
  ram[566]  = 255;
  ram[567]  = 255;
  ram[568]  = 255;
  ram[569]  = 255;
  ram[570]  = 255;
  ram[571]  = 255;
  ram[572]  = 255;
  ram[573]  = 255;
  ram[574]  = 255;
  ram[575]  = 255;
  ram[576]  = 255;
  ram[577]  = 255;
  ram[578]  = 255;
  ram[579]  = 255;
  ram[580]  = 255;
  ram[581]  = 255;
  ram[582]  = 255;
  ram[583]  = 255;
  ram[584]  = 255;
  ram[585]  = 255;
  ram[586]  = 255;
  ram[587]  = 255;
  ram[588]  = 255;
  ram[589]  = 255;
  ram[590]  = 255;
  ram[591]  = 255;
  ram[592]  = 255;
  ram[593]  = 255;
  ram[594]  = 255;
  ram[595]  = 255;
  ram[596]  = 255;
  ram[597]  = 255;
  ram[598]  = 255;
  ram[599]  = 255;
  ram[600]  = 255;
  ram[601]  = 255;
  ram[602]  = 255;
  ram[603]  = 255;
  ram[604]  = 255;
  ram[605]  = 255;
  ram[606]  = 255;
  ram[607]  = 255;
  ram[608]  = 255;
  ram[609]  = 255;
  ram[610]  = 255;
  ram[611]  = 255;
  ram[612]  = 255;
  ram[613]  = 255;
  ram[614]  = 255;
  ram[615]  = 255;
  ram[616]  = 255;
  ram[617]  = 255;
  ram[618]  = 255;
  ram[619]  = 255;
  ram[620]  = 255;
  ram[621]  = 255;
  ram[622]  = 255;
  ram[623]  = 255;
  ram[624]  = 255;
  ram[625]  = 255;
  ram[626]  = 255;
  ram[627]  = 255;
  ram[628]  = 255;
  ram[629]  = 255;
  ram[630]  = 255;
  ram[631]  = 255;
  ram[632]  = 255;
  ram[633]  = 255;
  ram[634]  = 255;
  ram[635]  = 255;
  ram[636]  = 255;
  ram[637]  = 255;
  ram[638]  = 255;
  ram[639]  = 255;
  ram[640]  = 255;
  ram[641]  = 255;
  ram[642]  = 255;
  ram[643]  = 255;
  ram[644]  = 255;
  ram[645]  = 255;
  ram[646]  = 255;
  ram[647]  = 255;
  ram[648]  = 255;
  ram[649]  = 255;
  ram[650]  = 255;
  ram[651]  = 255;
  ram[652]  = 255;
  ram[653]  = 255;
  ram[654]  = 255;
  ram[655]  = 255;
  ram[656]  = 255;
  ram[657]  = 255;
  ram[658]  = 255;
  ram[659]  = 255;
  ram[660]  = 255;
  ram[661]  = 255;
  ram[662]  = 255;
  ram[663]  = 255;
  ram[664]  = 255;
  ram[665]  = 255;
  ram[666]  = 255;
  ram[667]  = 255;
  ram[668]  = 255;
  ram[669]  = 255;
  ram[670]  = 255;
  ram[671]  = 255;
  ram[672]  = 255;
  ram[673]  = 255;
  ram[674]  = 255;
  ram[675]  = 255;
  ram[676]  = 255;
  ram[677]  = 255;
  ram[678]  = 255;
  ram[679]  = 255;
  ram[680]  = 255;
  ram[681]  = 255;
  ram[682]  = 255;
  ram[683]  = 255;
  ram[684]  = 255;
  ram[685]  = 255;
  ram[686]  = 255;
  ram[687]  = 255;
  ram[688]  = 255;
  ram[689]  = 255;
  ram[690]  = 255;
  ram[691]  = 255;
  ram[692]  = 255;
  ram[693]  = 255;
  ram[694]  = 255;
  ram[695]  = 255;
  ram[696]  = 255;
  ram[697]  = 255;
  ram[698]  = 255;
  ram[699]  = 255;
  ram[700]  = 255;
  ram[701]  = 255;
  ram[702]  = 255;
  ram[703]  = 255;
  ram[704]  = 255;
  ram[705]  = 255;
  ram[706]  = 255;
  ram[707]  = 255;
  ram[708]  = 255;
  ram[709]  = 255;
  ram[710]  = 255;
  ram[711]  = 255;
  ram[712]  = 255;
  ram[713]  = 255;
  ram[714]  = 255;
  ram[715]  = 255;
  ram[716]  = 255;
  ram[717]  = 255;
  ram[718]  = 255;
  ram[719]  = 255;
  ram[720]  = 255;
  ram[721]  = 255;
  ram[722]  = 255;
  ram[723]  = 255;
  ram[724]  = 255;
  ram[725]  = 255;
  ram[726]  = 255;
  ram[727]  = 255;
  ram[728]  = 255;
  ram[729]  = 255;
  ram[730]  = 255;
  ram[731]  = 255;
  ram[732]  = 255;
  ram[733]  = 255;
  ram[734]  = 255;
  ram[735]  = 255;
  ram[736]  = 255;
  ram[737]  = 255;
  ram[738]  = 255;
  ram[739]  = 255;
  ram[740]  = 255;
  ram[741]  = 255;
  ram[742]  = 255;
  ram[743]  = 255;
  ram[744]  = 255;
  ram[745]  = 255;
  ram[746]  = 255;
  ram[747]  = 255;
  ram[748]  = 255;
  ram[749]  = 255;
  ram[750]  = 255;
  ram[751]  = 255;
  ram[752]  = 255;
  ram[753]  = 255;
  ram[754]  = 255;
  ram[755]  = 255;
  ram[756]  = 255;
  ram[757]  = 255;
  ram[758]  = 255;
  ram[759]  = 255;
  ram[760]  = 255;
  ram[761]  = 255;
  ram[762]  = 255;
  ram[763]  = 255;
  ram[764]  = 255;
  ram[765]  = 255;
  ram[766]  = 255;
  ram[767]  = 255;
  ram[768]  = 255;
  ram[769]  = 255;
  ram[770]  = 255;
  ram[771]  = 255;
  ram[772]  = 255;
  ram[773]  = 255;
  ram[774]  = 255;
  ram[775]  = 255;
  ram[776]  = 255;
  ram[777]  = 255;
  ram[778]  = 255;
  ram[779]  = 255;
  ram[780]  = 255;
  ram[781]  = 255;
  ram[782]  = 255;
  ram[783]  = 255;
  ram[784]  = 255;
  ram[785]  = 255;
  ram[786]  = 255;
  ram[787]  = 255;
  ram[788]  = 255;
  ram[789]  = 255;
  ram[790]  = 255;
  ram[791]  = 255;
  ram[792]  = 255;
  ram[793]  = 255;
  ram[794]  = 255;
  ram[795]  = 255;
  ram[796]  = 255;
  ram[797]  = 255;
  ram[798]  = 255;
  ram[799]  = 255;
  ram[800]  = 255;
  ram[801]  = 255;
  ram[802]  = 255;
  ram[803]  = 255;
  ram[804]  = 255;
  ram[805]  = 255;
  ram[806]  = 255;
  ram[807]  = 255;
  ram[808]  = 255;
  ram[809]  = 255;
  ram[810]  = 255;
  ram[811]  = 255;
  ram[812]  = 255;
  ram[813]  = 255;
  ram[814]  = 255;
  ram[815]  = 255;
  ram[816]  = 255;
  ram[817]  = 255;
  ram[818]  = 255;
  ram[819]  = 255;
  ram[820]  = 255;
  ram[821]  = 255;
  ram[822]  = 181;
  ram[823]  = 122;
  ram[824]  = 71;
  ram[825]  = 71;
  ram[826]  = 71;
  ram[827]  = 71;
  ram[828]  = 137;
  ram[829]  = 181;
  ram[830]  = 236;
  ram[831]  = 255;
  ram[832]  = 255;
  ram[833]  = 255;
  ram[834]  = 255;
  ram[835]  = 255;
  ram[836]  = 255;
  ram[837]  = 255;
  ram[838]  = 255;
  ram[839]  = 221;
  ram[840]  = 137;
  ram[841]  = 137;
  ram[842]  = 167;
  ram[843]  = 255;
  ram[844]  = 255;
  ram[845]  = 255;
  ram[846]  = 255;
  ram[847]  = 255;
  ram[848]  = 255;
  ram[849]  = 255;
  ram[850]  = 255;
  ram[851]  = 255;
  ram[852]  = 255;
  ram[853]  = 167;
  ram[854]  = 137;
  ram[855]  = 167;
  ram[856]  = 255;
  ram[857]  = 255;
  ram[858]  = 255;
  ram[859]  = 255;
  ram[860]  = 255;
  ram[861]  = 255;
  ram[862]  = 255;
  ram[863]  = 255;
  ram[864]  = 255;
  ram[865]  = 255;
  ram[866]  = 255;
  ram[867]  = 255;
  ram[868]  = 255;
  ram[869]  = 255;
  ram[870]  = 255;
  ram[871]  = 255;
  ram[872]  = 255;
  ram[873]  = 255;
  ram[874]  = 255;
  ram[875]  = 255;
  ram[876]  = 255;
  ram[877]  = 255;
  ram[878]  = 255;
  ram[879]  = 255;
  ram[880]  = 255;
  ram[881]  = 255;
  ram[882]  = 255;
  ram[883]  = 255;
  ram[884]  = 255;
  ram[885]  = 255;
  ram[886]  = 255;
  ram[887]  = 255;
  ram[888]  = 255;
  ram[889]  = 255;
  ram[890]  = 255;
  ram[891]  = 255;
  ram[892]  = 255;
  ram[893]  = 255;
  ram[894]  = 255;
  ram[895]  = 255;
  ram[896]  = 255;
  ram[897]  = 255;
  ram[898]  = 255;
  ram[899]  = 255;
  ram[900]  = 137;
  ram[901]  = 17;
  ram[902]  = 0;
  ram[903]  = 0;
  ram[904]  = 0;
  ram[905]  = 0;
  ram[906]  = 0;
  ram[907]  = 0;
  ram[908]  = 0;
  ram[909]  = 0;
  ram[910]  = 137;
  ram[911]  = 255;
  ram[912]  = 255;
  ram[913]  = 255;
  ram[914]  = 255;
  ram[915]  = 255;
  ram[916]  = 255;
  ram[917]  = 255;
  ram[918]  = 255;
  ram[919]  = 122;
  ram[920]  = 0;
  ram[921]  = 0;
  ram[922]  = 17;
  ram[923]  = 236;
  ram[924]  = 255;
  ram[925]  = 255;
  ram[926]  = 255;
  ram[927]  = 255;
  ram[928]  = 255;
  ram[929]  = 255;
  ram[930]  = 255;
  ram[931]  = 255;
  ram[932]  = 255;
  ram[933]  = 71;
  ram[934]  = 0;
  ram[935]  = 71;
  ram[936]  = 255;
  ram[937]  = 255;
  ram[938]  = 255;
  ram[939]  = 255;
  ram[940]  = 255;
  ram[941]  = 255;
  ram[942]  = 255;
  ram[943]  = 255;
  ram[944]  = 255;
  ram[945]  = 255;
  ram[946]  = 255;
  ram[947]  = 255;
  ram[948]  = 255;
  ram[949]  = 255;
  ram[950]  = 255;
  ram[951]  = 255;
  ram[952]  = 255;
  ram[953]  = 255;
  ram[954]  = 255;
  ram[955]  = 255;
  ram[956]  = 255;
  ram[957]  = 255;
  ram[958]  = 255;
  ram[959]  = 255;
  ram[960]  = 255;
  ram[961]  = 255;
  ram[962]  = 255;
  ram[963]  = 255;
  ram[964]  = 255;
  ram[965]  = 255;
  ram[966]  = 255;
  ram[967]  = 255;
  ram[968]  = 255;
  ram[969]  = 255;
  ram[970]  = 255;
  ram[971]  = 255;
  ram[972]  = 255;
  ram[973]  = 255;
  ram[974]  = 255;
  ram[975]  = 255;
  ram[976]  = 255;
  ram[977]  = 255;
  ram[978]  = 236;
  ram[979]  = 52;
  ram[980]  = 0;
  ram[981]  = 0;
  ram[982]  = 0;
  ram[983]  = 35;
  ram[984]  = 71;
  ram[985]  = 122;
  ram[986]  = 105;
  ram[987]  = 71;
  ram[988]  = 17;
  ram[989]  = 0;
  ram[990]  = 137;
  ram[991]  = 255;
  ram[992]  = 255;
  ram[993]  = 255;
  ram[994]  = 255;
  ram[995]  = 255;
  ram[996]  = 255;
  ram[997]  = 255;
  ram[998]  = 255;
  ram[999]  = 35;
  ram[1000]  = 0;
  ram[1001]  = 0;
  ram[1002]  = 0;
  ram[1003]  = 167;
  ram[1004]  = 255;
  ram[1005]  = 255;
  ram[1006]  = 255;
  ram[1007]  = 255;
  ram[1008]  = 255;
  ram[1009]  = 255;
  ram[1010]  = 255;
  ram[1011]  = 255;
  ram[1012]  = 255;
  ram[1013]  = 71;
  ram[1014]  = 0;
  ram[1015]  = 71;
  ram[1016]  = 255;
  ram[1017]  = 255;
  ram[1018]  = 255;
  ram[1019]  = 255;
  ram[1020]  = 255;
  ram[1021]  = 255;
  ram[1022]  = 255;
  ram[1023]  = 255;
  ram[1024]  = 255;
  ram[1025]  = 255;
  ram[1026]  = 255;
  ram[1027]  = 255;
  ram[1028]  = 255;
  ram[1029]  = 255;
  ram[1030]  = 255;
  ram[1031]  = 255;
  ram[1032]  = 255;
  ram[1033]  = 255;
  ram[1034]  = 255;
  ram[1035]  = 255;
  ram[1036]  = 255;
  ram[1037]  = 255;
  ram[1038]  = 255;
  ram[1039]  = 255;
  ram[1040]  = 255;
  ram[1041]  = 255;
  ram[1042]  = 255;
  ram[1043]  = 255;
  ram[1044]  = 255;
  ram[1045]  = 255;
  ram[1046]  = 255;
  ram[1047]  = 255;
  ram[1048]  = 255;
  ram[1049]  = 255;
  ram[1050]  = 255;
  ram[1051]  = 255;
  ram[1052]  = 255;
  ram[1053]  = 255;
  ram[1054]  = 255;
  ram[1055]  = 255;
  ram[1056]  = 255;
  ram[1057]  = 236;
  ram[1058]  = 52;
  ram[1059]  = 0;
  ram[1060]  = 0;
  ram[1061]  = 52;
  ram[1062]  = 195;
  ram[1063]  = 255;
  ram[1064]  = 255;
  ram[1065]  = 255;
  ram[1066]  = 255;
  ram[1067]  = 255;
  ram[1068]  = 255;
  ram[1069]  = 181;
  ram[1070]  = 181;
  ram[1071]  = 255;
  ram[1072]  = 255;
  ram[1073]  = 255;
  ram[1074]  = 255;
  ram[1075]  = 255;
  ram[1076]  = 255;
  ram[1077]  = 255;
  ram[1078]  = 181;
  ram[1079]  = 0;
  ram[1080]  = 0;
  ram[1081]  = 52;
  ram[1082]  = 0;
  ram[1083]  = 52;
  ram[1084]  = 255;
  ram[1085]  = 255;
  ram[1086]  = 255;
  ram[1087]  = 255;
  ram[1088]  = 255;
  ram[1089]  = 255;
  ram[1090]  = 255;
  ram[1091]  = 255;
  ram[1092]  = 255;
  ram[1093]  = 71;
  ram[1094]  = 0;
  ram[1095]  = 71;
  ram[1096]  = 255;
  ram[1097]  = 255;
  ram[1098]  = 255;
  ram[1099]  = 255;
  ram[1100]  = 255;
  ram[1101]  = 255;
  ram[1102]  = 255;
  ram[1103]  = 255;
  ram[1104]  = 255;
  ram[1105]  = 255;
  ram[1106]  = 255;
  ram[1107]  = 255;
  ram[1108]  = 255;
  ram[1109]  = 255;
  ram[1110]  = 255;
  ram[1111]  = 255;
  ram[1112]  = 255;
  ram[1113]  = 255;
  ram[1114]  = 255;
  ram[1115]  = 255;
  ram[1116]  = 255;
  ram[1117]  = 255;
  ram[1118]  = 255;
  ram[1119]  = 255;
  ram[1120]  = 255;
  ram[1121]  = 255;
  ram[1122]  = 255;
  ram[1123]  = 255;
  ram[1124]  = 255;
  ram[1125]  = 255;
  ram[1126]  = 255;
  ram[1127]  = 255;
  ram[1128]  = 255;
  ram[1129]  = 255;
  ram[1130]  = 255;
  ram[1131]  = 255;
  ram[1132]  = 255;
  ram[1133]  = 255;
  ram[1134]  = 255;
  ram[1135]  = 255;
  ram[1136]  = 255;
  ram[1137]  = 71;
  ram[1138]  = 0;
  ram[1139]  = 0;
  ram[1140]  = 105;
  ram[1141]  = 255;
  ram[1142]  = 255;
  ram[1143]  = 255;
  ram[1144]  = 255;
  ram[1145]  = 255;
  ram[1146]  = 255;
  ram[1147]  = 255;
  ram[1148]  = 255;
  ram[1149]  = 255;
  ram[1150]  = 255;
  ram[1151]  = 255;
  ram[1152]  = 255;
  ram[1153]  = 255;
  ram[1154]  = 255;
  ram[1155]  = 255;
  ram[1156]  = 255;
  ram[1157]  = 255;
  ram[1158]  = 105;
  ram[1159]  = 0;
  ram[1160]  = 35;
  ram[1161]  = 152;
  ram[1162]  = 0;
  ram[1163]  = 0;
  ram[1164]  = 221;
  ram[1165]  = 255;
  ram[1166]  = 255;
  ram[1167]  = 255;
  ram[1168]  = 255;
  ram[1169]  = 255;
  ram[1170]  = 255;
  ram[1171]  = 255;
  ram[1172]  = 255;
  ram[1173]  = 71;
  ram[1174]  = 0;
  ram[1175]  = 71;
  ram[1176]  = 255;
  ram[1177]  = 255;
  ram[1178]  = 255;
  ram[1179]  = 255;
  ram[1180]  = 255;
  ram[1181]  = 255;
  ram[1182]  = 255;
  ram[1183]  = 255;
  ram[1184]  = 255;
  ram[1185]  = 255;
  ram[1186]  = 255;
  ram[1187]  = 255;
  ram[1188]  = 255;
  ram[1189]  = 255;
  ram[1190]  = 255;
  ram[1191]  = 255;
  ram[1192]  = 255;
  ram[1193]  = 255;
  ram[1194]  = 255;
  ram[1195]  = 255;
  ram[1196]  = 255;
  ram[1197]  = 255;
  ram[1198]  = 255;
  ram[1199]  = 255;
  ram[1200]  = 255;
  ram[1201]  = 255;
  ram[1202]  = 255;
  ram[1203]  = 255;
  ram[1204]  = 255;
  ram[1205]  = 255;
  ram[1206]  = 255;
  ram[1207]  = 255;
  ram[1208]  = 255;
  ram[1209]  = 255;
  ram[1210]  = 255;
  ram[1211]  = 255;
  ram[1212]  = 255;
  ram[1213]  = 255;
  ram[1214]  = 255;
  ram[1215]  = 255;
  ram[1216]  = 167;
  ram[1217]  = 0;
  ram[1218]  = 0;
  ram[1219]  = 71;
  ram[1220]  = 255;
  ram[1221]  = 255;
  ram[1222]  = 255;
  ram[1223]  = 255;
  ram[1224]  = 255;
  ram[1225]  = 255;
  ram[1226]  = 255;
  ram[1227]  = 255;
  ram[1228]  = 255;
  ram[1229]  = 255;
  ram[1230]  = 255;
  ram[1231]  = 255;
  ram[1232]  = 255;
  ram[1233]  = 255;
  ram[1234]  = 255;
  ram[1235]  = 255;
  ram[1236]  = 255;
  ram[1237]  = 236;
  ram[1238]  = 0;
  ram[1239]  = 0;
  ram[1240]  = 137;
  ram[1241]  = 221;
  ram[1242]  = 0;
  ram[1243]  = 0;
  ram[1244]  = 122;
  ram[1245]  = 255;
  ram[1246]  = 255;
  ram[1247]  = 255;
  ram[1248]  = 255;
  ram[1249]  = 255;
  ram[1250]  = 255;
  ram[1251]  = 255;
  ram[1252]  = 255;
  ram[1253]  = 71;
  ram[1254]  = 0;
  ram[1255]  = 71;
  ram[1256]  = 255;
  ram[1257]  = 255;
  ram[1258]  = 255;
  ram[1259]  = 255;
  ram[1260]  = 255;
  ram[1261]  = 255;
  ram[1262]  = 255;
  ram[1263]  = 255;
  ram[1264]  = 255;
  ram[1265]  = 255;
  ram[1266]  = 255;
  ram[1267]  = 255;
  ram[1268]  = 255;
  ram[1269]  = 255;
  ram[1270]  = 255;
  ram[1271]  = 255;
  ram[1272]  = 255;
  ram[1273]  = 255;
  ram[1274]  = 255;
  ram[1275]  = 255;
  ram[1276]  = 255;
  ram[1277]  = 255;
  ram[1278]  = 255;
  ram[1279]  = 255;
  ram[1280]  = 255;
  ram[1281]  = 255;
  ram[1282]  = 255;
  ram[1283]  = 255;
  ram[1284]  = 255;
  ram[1285]  = 255;
  ram[1286]  = 255;
  ram[1287]  = 255;
  ram[1288]  = 255;
  ram[1289]  = 255;
  ram[1290]  = 255;
  ram[1291]  = 255;
  ram[1292]  = 255;
  ram[1293]  = 255;
  ram[1294]  = 255;
  ram[1295]  = 255;
  ram[1296]  = 35;
  ram[1297]  = 0;
  ram[1298]  = 0;
  ram[1299]  = 221;
  ram[1300]  = 255;
  ram[1301]  = 255;
  ram[1302]  = 255;
  ram[1303]  = 255;
  ram[1304]  = 255;
  ram[1305]  = 255;
  ram[1306]  = 255;
  ram[1307]  = 255;
  ram[1308]  = 255;
  ram[1309]  = 255;
  ram[1310]  = 255;
  ram[1311]  = 255;
  ram[1312]  = 255;
  ram[1313]  = 255;
  ram[1314]  = 255;
  ram[1315]  = 255;
  ram[1316]  = 255;
  ram[1317]  = 152;
  ram[1318]  = 0;
  ram[1319]  = 0;
  ram[1320]  = 221;
  ram[1321]  = 255;
  ram[1322]  = 52;
  ram[1323]  = 0;
  ram[1324]  = 35;
  ram[1325]  = 255;
  ram[1326]  = 255;
  ram[1327]  = 255;
  ram[1328]  = 255;
  ram[1329]  = 255;
  ram[1330]  = 255;
  ram[1331]  = 255;
  ram[1332]  = 255;
  ram[1333]  = 71;
  ram[1334]  = 0;
  ram[1335]  = 71;
  ram[1336]  = 255;
  ram[1337]  = 255;
  ram[1338]  = 255;
  ram[1339]  = 255;
  ram[1340]  = 255;
  ram[1341]  = 255;
  ram[1342]  = 255;
  ram[1343]  = 255;
  ram[1344]  = 255;
  ram[1345]  = 255;
  ram[1346]  = 255;
  ram[1347]  = 255;
  ram[1348]  = 255;
  ram[1349]  = 255;
  ram[1350]  = 255;
  ram[1351]  = 255;
  ram[1352]  = 255;
  ram[1353]  = 255;
  ram[1354]  = 255;
  ram[1355]  = 255;
  ram[1356]  = 255;
  ram[1357]  = 255;
  ram[1358]  = 255;
  ram[1359]  = 255;
  ram[1360]  = 255;
  ram[1361]  = 255;
  ram[1362]  = 255;
  ram[1363]  = 255;
  ram[1364]  = 255;
  ram[1365]  = 255;
  ram[1366]  = 255;
  ram[1367]  = 255;
  ram[1368]  = 255;
  ram[1369]  = 255;
  ram[1370]  = 255;
  ram[1371]  = 255;
  ram[1372]  = 255;
  ram[1373]  = 255;
  ram[1374]  = 255;
  ram[1375]  = 208;
  ram[1376]  = 0;
  ram[1377]  = 0;
  ram[1378]  = 105;
  ram[1379]  = 255;
  ram[1380]  = 255;
  ram[1381]  = 255;
  ram[1382]  = 255;
  ram[1383]  = 255;
  ram[1384]  = 255;
  ram[1385]  = 255;
  ram[1386]  = 255;
  ram[1387]  = 255;
  ram[1388]  = 255;
  ram[1389]  = 255;
  ram[1390]  = 255;
  ram[1391]  = 255;
  ram[1392]  = 255;
  ram[1393]  = 255;
  ram[1394]  = 255;
  ram[1395]  = 255;
  ram[1396]  = 255;
  ram[1397]  = 52;
  ram[1398]  = 0;
  ram[1399]  = 52;
  ram[1400]  = 255;
  ram[1401]  = 255;
  ram[1402]  = 167;
  ram[1403]  = 0;
  ram[1404]  = 0;
  ram[1405]  = 181;
  ram[1406]  = 255;
  ram[1407]  = 255;
  ram[1408]  = 255;
  ram[1409]  = 255;
  ram[1410]  = 255;
  ram[1411]  = 255;
  ram[1412]  = 255;
  ram[1413]  = 71;
  ram[1414]  = 0;
  ram[1415]  = 71;
  ram[1416]  = 255;
  ram[1417]  = 255;
  ram[1418]  = 255;
  ram[1419]  = 255;
  ram[1420]  = 255;
  ram[1421]  = 255;
  ram[1422]  = 255;
  ram[1423]  = 255;
  ram[1424]  = 255;
  ram[1425]  = 255;
  ram[1426]  = 255;
  ram[1427]  = 255;
  ram[1428]  = 255;
  ram[1429]  = 255;
  ram[1430]  = 255;
  ram[1431]  = 255;
  ram[1432]  = 255;
  ram[1433]  = 255;
  ram[1434]  = 255;
  ram[1435]  = 255;
  ram[1436]  = 255;
  ram[1437]  = 255;
  ram[1438]  = 255;
  ram[1439]  = 255;
  ram[1440]  = 255;
  ram[1441]  = 255;
  ram[1442]  = 255;
  ram[1443]  = 255;
  ram[1444]  = 255;
  ram[1445]  = 255;
  ram[1446]  = 255;
  ram[1447]  = 255;
  ram[1448]  = 255;
  ram[1449]  = 255;
  ram[1450]  = 255;
  ram[1451]  = 255;
  ram[1452]  = 255;
  ram[1453]  = 255;
  ram[1454]  = 255;
  ram[1455]  = 152;
  ram[1456]  = 0;
  ram[1457]  = 0;
  ram[1458]  = 167;
  ram[1459]  = 255;
  ram[1460]  = 255;
  ram[1461]  = 255;
  ram[1462]  = 255;
  ram[1463]  = 255;
  ram[1464]  = 255;
  ram[1465]  = 255;
  ram[1466]  = 255;
  ram[1467]  = 255;
  ram[1468]  = 255;
  ram[1469]  = 255;
  ram[1470]  = 255;
  ram[1471]  = 255;
  ram[1472]  = 255;
  ram[1473]  = 255;
  ram[1474]  = 255;
  ram[1475]  = 255;
  ram[1476]  = 208;
  ram[1477]  = 0;
  ram[1478]  = 0;
  ram[1479]  = 152;
  ram[1480]  = 255;
  ram[1481]  = 255;
  ram[1482]  = 236;
  ram[1483]  = 0;
  ram[1484]  = 0;
  ram[1485]  = 87;
  ram[1486]  = 255;
  ram[1487]  = 255;
  ram[1488]  = 255;
  ram[1489]  = 255;
  ram[1490]  = 255;
  ram[1491]  = 255;
  ram[1492]  = 255;
  ram[1493]  = 71;
  ram[1494]  = 0;
  ram[1495]  = 71;
  ram[1496]  = 255;
  ram[1497]  = 255;
  ram[1498]  = 255;
  ram[1499]  = 255;
  ram[1500]  = 255;
  ram[1501]  = 255;
  ram[1502]  = 255;
  ram[1503]  = 255;
  ram[1504]  = 255;
  ram[1505]  = 255;
  ram[1506]  = 255;
  ram[1507]  = 255;
  ram[1508]  = 255;
  ram[1509]  = 255;
  ram[1510]  = 255;
  ram[1511]  = 255;
  ram[1512]  = 255;
  ram[1513]  = 255;
  ram[1514]  = 255;
  ram[1515]  = 255;
  ram[1516]  = 255;
  ram[1517]  = 255;
  ram[1518]  = 255;
  ram[1519]  = 255;
  ram[1520]  = 255;
  ram[1521]  = 255;
  ram[1522]  = 255;
  ram[1523]  = 255;
  ram[1524]  = 255;
  ram[1525]  = 255;
  ram[1526]  = 255;
  ram[1527]  = 255;
  ram[1528]  = 255;
  ram[1529]  = 255;
  ram[1530]  = 255;
  ram[1531]  = 255;
  ram[1532]  = 255;
  ram[1533]  = 255;
  ram[1534]  = 255;
  ram[1535]  = 122;
  ram[1536]  = 0;
  ram[1537]  = 0;
  ram[1538]  = 195;
  ram[1539]  = 255;
  ram[1540]  = 255;
  ram[1541]  = 255;
  ram[1542]  = 255;
  ram[1543]  = 255;
  ram[1544]  = 255;
  ram[1545]  = 255;
  ram[1546]  = 255;
  ram[1547]  = 255;
  ram[1548]  = 255;
  ram[1549]  = 255;
  ram[1550]  = 255;
  ram[1551]  = 255;
  ram[1552]  = 255;
  ram[1553]  = 255;
  ram[1554]  = 255;
  ram[1555]  = 255;
  ram[1556]  = 122;
  ram[1557]  = 0;
  ram[1558]  = 0;
  ram[1559]  = 236;
  ram[1560]  = 255;
  ram[1561]  = 255;
  ram[1562]  = 255;
  ram[1563]  = 87;
  ram[1564]  = 0;
  ram[1565]  = 0;
  ram[1566]  = 236;
  ram[1567]  = 255;
  ram[1568]  = 255;
  ram[1569]  = 255;
  ram[1570]  = 255;
  ram[1571]  = 255;
  ram[1572]  = 255;
  ram[1573]  = 71;
  ram[1574]  = 0;
  ram[1575]  = 71;
  ram[1576]  = 255;
  ram[1577]  = 255;
  ram[1578]  = 255;
  ram[1579]  = 255;
  ram[1580]  = 255;
  ram[1581]  = 255;
  ram[1582]  = 255;
  ram[1583]  = 255;
  ram[1584]  = 255;
  ram[1585]  = 255;
  ram[1586]  = 255;
  ram[1587]  = 255;
  ram[1588]  = 255;
  ram[1589]  = 255;
  ram[1590]  = 255;
  ram[1591]  = 255;
  ram[1592]  = 255;
  ram[1593]  = 255;
  ram[1594]  = 255;
  ram[1595]  = 255;
  ram[1596]  = 255;
  ram[1597]  = 255;
  ram[1598]  = 255;
  ram[1599]  = 255;
  ram[1600]  = 255;
  ram[1601]  = 255;
  ram[1602]  = 255;
  ram[1603]  = 255;
  ram[1604]  = 255;
  ram[1605]  = 255;
  ram[1606]  = 255;
  ram[1607]  = 255;
  ram[1608]  = 255;
  ram[1609]  = 255;
  ram[1610]  = 255;
  ram[1611]  = 255;
  ram[1612]  = 255;
  ram[1613]  = 255;
  ram[1614]  = 255;
  ram[1615]  = 71;
  ram[1616]  = 0;
  ram[1617]  = 0;
  ram[1618]  = 255;
  ram[1619]  = 255;
  ram[1620]  = 255;
  ram[1621]  = 255;
  ram[1622]  = 255;
  ram[1623]  = 255;
  ram[1624]  = 255;
  ram[1625]  = 255;
  ram[1626]  = 255;
  ram[1627]  = 255;
  ram[1628]  = 255;
  ram[1629]  = 255;
  ram[1630]  = 255;
  ram[1631]  = 255;
  ram[1632]  = 255;
  ram[1633]  = 255;
  ram[1634]  = 255;
  ram[1635]  = 255;
  ram[1636]  = 17;
  ram[1637]  = 0;
  ram[1638]  = 87;
  ram[1639]  = 255;
  ram[1640]  = 255;
  ram[1641]  = 255;
  ram[1642]  = 255;
  ram[1643]  = 181;
  ram[1644]  = 0;
  ram[1645]  = 0;
  ram[1646]  = 152;
  ram[1647]  = 255;
  ram[1648]  = 255;
  ram[1649]  = 255;
  ram[1650]  = 255;
  ram[1651]  = 255;
  ram[1652]  = 255;
  ram[1653]  = 71;
  ram[1654]  = 0;
  ram[1655]  = 71;
  ram[1656]  = 255;
  ram[1657]  = 255;
  ram[1658]  = 255;
  ram[1659]  = 255;
  ram[1660]  = 255;
  ram[1661]  = 255;
  ram[1662]  = 255;
  ram[1663]  = 255;
  ram[1664]  = 255;
  ram[1665]  = 255;
  ram[1666]  = 255;
  ram[1667]  = 255;
  ram[1668]  = 255;
  ram[1669]  = 255;
  ram[1670]  = 255;
  ram[1671]  = 255;
  ram[1672]  = 255;
  ram[1673]  = 255;
  ram[1674]  = 255;
  ram[1675]  = 255;
  ram[1676]  = 255;
  ram[1677]  = 255;
  ram[1678]  = 255;
  ram[1679]  = 255;
  ram[1680]  = 255;
  ram[1681]  = 255;
  ram[1682]  = 255;
  ram[1683]  = 255;
  ram[1684]  = 255;
  ram[1685]  = 255;
  ram[1686]  = 255;
  ram[1687]  = 255;
  ram[1688]  = 255;
  ram[1689]  = 255;
  ram[1690]  = 255;
  ram[1691]  = 255;
  ram[1692]  = 255;
  ram[1693]  = 255;
  ram[1694]  = 255;
  ram[1695]  = 71;
  ram[1696]  = 0;
  ram[1697]  = 0;
  ram[1698]  = 255;
  ram[1699]  = 255;
  ram[1700]  = 255;
  ram[1701]  = 255;
  ram[1702]  = 255;
  ram[1703]  = 255;
  ram[1704]  = 255;
  ram[1705]  = 255;
  ram[1706]  = 255;
  ram[1707]  = 255;
  ram[1708]  = 255;
  ram[1709]  = 255;
  ram[1710]  = 255;
  ram[1711]  = 255;
  ram[1712]  = 255;
  ram[1713]  = 255;
  ram[1714]  = 255;
  ram[1715]  = 167;
  ram[1716]  = 0;
  ram[1717]  = 0;
  ram[1718]  = 167;
  ram[1719]  = 255;
  ram[1720]  = 255;
  ram[1721]  = 255;
  ram[1722]  = 255;
  ram[1723]  = 255;
  ram[1724]  = 17;
  ram[1725]  = 0;
  ram[1726]  = 52;
  ram[1727]  = 255;
  ram[1728]  = 255;
  ram[1729]  = 255;
  ram[1730]  = 255;
  ram[1731]  = 255;
  ram[1732]  = 255;
  ram[1733]  = 71;
  ram[1734]  = 0;
  ram[1735]  = 71;
  ram[1736]  = 255;
  ram[1737]  = 255;
  ram[1738]  = 255;
  ram[1739]  = 255;
  ram[1740]  = 255;
  ram[1741]  = 255;
  ram[1742]  = 255;
  ram[1743]  = 255;
  ram[1744]  = 255;
  ram[1745]  = 255;
  ram[1746]  = 255;
  ram[1747]  = 255;
  ram[1748]  = 255;
  ram[1749]  = 255;
  ram[1750]  = 255;
  ram[1751]  = 255;
  ram[1752]  = 255;
  ram[1753]  = 255;
  ram[1754]  = 255;
  ram[1755]  = 255;
  ram[1756]  = 255;
  ram[1757]  = 255;
  ram[1758]  = 255;
  ram[1759]  = 255;
  ram[1760]  = 255;
  ram[1761]  = 255;
  ram[1762]  = 255;
  ram[1763]  = 255;
  ram[1764]  = 255;
  ram[1765]  = 255;
  ram[1766]  = 255;
  ram[1767]  = 255;
  ram[1768]  = 255;
  ram[1769]  = 255;
  ram[1770]  = 255;
  ram[1771]  = 255;
  ram[1772]  = 255;
  ram[1773]  = 255;
  ram[1774]  = 255;
  ram[1775]  = 105;
  ram[1776]  = 0;
  ram[1777]  = 0;
  ram[1778]  = 195;
  ram[1779]  = 255;
  ram[1780]  = 255;
  ram[1781]  = 255;
  ram[1782]  = 255;
  ram[1783]  = 255;
  ram[1784]  = 255;
  ram[1785]  = 255;
  ram[1786]  = 255;
  ram[1787]  = 255;
  ram[1788]  = 255;
  ram[1789]  = 255;
  ram[1790]  = 255;
  ram[1791]  = 255;
  ram[1792]  = 255;
  ram[1793]  = 255;
  ram[1794]  = 255;
  ram[1795]  = 87;
  ram[1796]  = 0;
  ram[1797]  = 17;
  ram[1798]  = 255;
  ram[1799]  = 255;
  ram[1800]  = 255;
  ram[1801]  = 255;
  ram[1802]  = 255;
  ram[1803]  = 255;
  ram[1804]  = 105;
  ram[1805]  = 0;
  ram[1806]  = 0;
  ram[1807]  = 208;
  ram[1808]  = 255;
  ram[1809]  = 255;
  ram[1810]  = 255;
  ram[1811]  = 255;
  ram[1812]  = 255;
  ram[1813]  = 71;
  ram[1814]  = 0;
  ram[1815]  = 71;
  ram[1816]  = 255;
  ram[1817]  = 255;
  ram[1818]  = 255;
  ram[1819]  = 255;
  ram[1820]  = 255;
  ram[1821]  = 255;
  ram[1822]  = 255;
  ram[1823]  = 255;
  ram[1824]  = 255;
  ram[1825]  = 255;
  ram[1826]  = 255;
  ram[1827]  = 255;
  ram[1828]  = 255;
  ram[1829]  = 255;
  ram[1830]  = 255;
  ram[1831]  = 255;
  ram[1832]  = 255;
  ram[1833]  = 255;
  ram[1834]  = 255;
  ram[1835]  = 255;
  ram[1836]  = 255;
  ram[1837]  = 255;
  ram[1838]  = 255;
  ram[1839]  = 255;
  ram[1840]  = 255;
  ram[1841]  = 255;
  ram[1842]  = 255;
  ram[1843]  = 255;
  ram[1844]  = 255;
  ram[1845]  = 255;
  ram[1846]  = 255;
  ram[1847]  = 255;
  ram[1848]  = 255;
  ram[1849]  = 255;
  ram[1850]  = 255;
  ram[1851]  = 255;
  ram[1852]  = 255;
  ram[1853]  = 255;
  ram[1854]  = 255;
  ram[1855]  = 137;
  ram[1856]  = 0;
  ram[1857]  = 0;
  ram[1858]  = 167;
  ram[1859]  = 255;
  ram[1860]  = 255;
  ram[1861]  = 255;
  ram[1862]  = 255;
  ram[1863]  = 255;
  ram[1864]  = 255;
  ram[1865]  = 255;
  ram[1866]  = 255;
  ram[1867]  = 255;
  ram[1868]  = 255;
  ram[1869]  = 255;
  ram[1870]  = 255;
  ram[1871]  = 255;
  ram[1872]  = 255;
  ram[1873]  = 255;
  ram[1874]  = 221;
  ram[1875]  = 0;
  ram[1876]  = 0;
  ram[1877]  = 0;
  ram[1878]  = 0;
  ram[1879]  = 0;
  ram[1880]  = 0;
  ram[1881]  = 0;
  ram[1882]  = 0;
  ram[1883]  = 0;
  ram[1884]  = 0;
  ram[1885]  = 0;
  ram[1886]  = 0;
  ram[1887]  = 105;
  ram[1888]  = 255;
  ram[1889]  = 255;
  ram[1890]  = 255;
  ram[1891]  = 255;
  ram[1892]  = 255;
  ram[1893]  = 71;
  ram[1894]  = 0;
  ram[1895]  = 71;
  ram[1896]  = 255;
  ram[1897]  = 255;
  ram[1898]  = 255;
  ram[1899]  = 255;
  ram[1900]  = 255;
  ram[1901]  = 255;
  ram[1902]  = 255;
  ram[1903]  = 255;
  ram[1904]  = 255;
  ram[1905]  = 255;
  ram[1906]  = 255;
  ram[1907]  = 255;
  ram[1908]  = 255;
  ram[1909]  = 255;
  ram[1910]  = 255;
  ram[1911]  = 255;
  ram[1912]  = 255;
  ram[1913]  = 255;
  ram[1914]  = 255;
  ram[1915]  = 255;
  ram[1916]  = 255;
  ram[1917]  = 255;
  ram[1918]  = 255;
  ram[1919]  = 255;
  ram[1920]  = 255;
  ram[1921]  = 255;
  ram[1922]  = 255;
  ram[1923]  = 255;
  ram[1924]  = 255;
  ram[1925]  = 255;
  ram[1926]  = 255;
  ram[1927]  = 255;
  ram[1928]  = 255;
  ram[1929]  = 255;
  ram[1930]  = 255;
  ram[1931]  = 255;
  ram[1932]  = 255;
  ram[1933]  = 255;
  ram[1934]  = 255;
  ram[1935]  = 181;
  ram[1936]  = 0;
  ram[1937]  = 0;
  ram[1938]  = 105;
  ram[1939]  = 255;
  ram[1940]  = 255;
  ram[1941]  = 255;
  ram[1942]  = 255;
  ram[1943]  = 255;
  ram[1944]  = 255;
  ram[1945]  = 255;
  ram[1946]  = 255;
  ram[1947]  = 255;
  ram[1948]  = 255;
  ram[1949]  = 255;
  ram[1950]  = 255;
  ram[1951]  = 255;
  ram[1952]  = 255;
  ram[1953]  = 255;
  ram[1954]  = 152;
  ram[1955]  = 0;
  ram[1956]  = 0;
  ram[1957]  = 0;
  ram[1958]  = 0;
  ram[1959]  = 0;
  ram[1960]  = 0;
  ram[1961]  = 0;
  ram[1962]  = 0;
  ram[1963]  = 0;
  ram[1964]  = 0;
  ram[1965]  = 0;
  ram[1966]  = 0;
  ram[1967]  = 17;
  ram[1968]  = 255;
  ram[1969]  = 255;
  ram[1970]  = 255;
  ram[1971]  = 255;
  ram[1972]  = 255;
  ram[1973]  = 71;
  ram[1974]  = 0;
  ram[1975]  = 71;
  ram[1976]  = 255;
  ram[1977]  = 255;
  ram[1978]  = 255;
  ram[1979]  = 255;
  ram[1980]  = 255;
  ram[1981]  = 255;
  ram[1982]  = 255;
  ram[1983]  = 255;
  ram[1984]  = 255;
  ram[1985]  = 255;
  ram[1986]  = 255;
  ram[1987]  = 255;
  ram[1988]  = 255;
  ram[1989]  = 255;
  ram[1990]  = 255;
  ram[1991]  = 255;
  ram[1992]  = 255;
  ram[1993]  = 255;
  ram[1994]  = 255;
  ram[1995]  = 255;
  ram[1996]  = 255;
  ram[1997]  = 255;
  ram[1998]  = 255;
  ram[1999]  = 255;
  ram[2000]  = 255;
  ram[2001]  = 255;
  ram[2002]  = 255;
  ram[2003]  = 255;
  ram[2004]  = 255;
  ram[2005]  = 255;
  ram[2006]  = 255;
  ram[2007]  = 255;
  ram[2008]  = 255;
  ram[2009]  = 255;
  ram[2010]  = 255;
  ram[2011]  = 255;
  ram[2012]  = 255;
  ram[2013]  = 255;
  ram[2014]  = 255;
  ram[2015]  = 255;
  ram[2016]  = 17;
  ram[2017]  = 0;
  ram[2018]  = 0;
  ram[2019]  = 221;
  ram[2020]  = 255;
  ram[2021]  = 255;
  ram[2022]  = 255;
  ram[2023]  = 255;
  ram[2024]  = 255;
  ram[2025]  = 255;
  ram[2026]  = 255;
  ram[2027]  = 255;
  ram[2028]  = 255;
  ram[2029]  = 255;
  ram[2030]  = 255;
  ram[2031]  = 255;
  ram[2032]  = 255;
  ram[2033]  = 255;
  ram[2034]  = 35;
  ram[2035]  = 0;
  ram[2036]  = 35;
  ram[2037]  = 137;
  ram[2038]  = 137;
  ram[2039]  = 137;
  ram[2040]  = 137;
  ram[2041]  = 137;
  ram[2042]  = 137;
  ram[2043]  = 137;
  ram[2044]  = 137;
  ram[2045]  = 71;
  ram[2046]  = 0;
  ram[2047]  = 0;
  ram[2048]  = 167;
  ram[2049]  = 255;
  ram[2050]  = 255;
  ram[2051]  = 255;
  ram[2052]  = 255;
  ram[2053]  = 71;
  ram[2054]  = 0;
  ram[2055]  = 71;
  ram[2056]  = 255;
  ram[2057]  = 255;
  ram[2058]  = 255;
  ram[2059]  = 255;
  ram[2060]  = 255;
  ram[2061]  = 255;
  ram[2062]  = 255;
  ram[2063]  = 255;
  ram[2064]  = 255;
  ram[2065]  = 255;
  ram[2066]  = 255;
  ram[2067]  = 255;
  ram[2068]  = 255;
  ram[2069]  = 255;
  ram[2070]  = 255;
  ram[2071]  = 255;
  ram[2072]  = 255;
  ram[2073]  = 255;
  ram[2074]  = 255;
  ram[2075]  = 255;
  ram[2076]  = 255;
  ram[2077]  = 255;
  ram[2078]  = 255;
  ram[2079]  = 255;
  ram[2080]  = 255;
  ram[2081]  = 255;
  ram[2082]  = 255;
  ram[2083]  = 255;
  ram[2084]  = 255;
  ram[2085]  = 255;
  ram[2086]  = 255;
  ram[2087]  = 255;
  ram[2088]  = 255;
  ram[2089]  = 255;
  ram[2090]  = 255;
  ram[2091]  = 255;
  ram[2092]  = 255;
  ram[2093]  = 255;
  ram[2094]  = 255;
  ram[2095]  = 255;
  ram[2096]  = 137;
  ram[2097]  = 0;
  ram[2098]  = 0;
  ram[2099]  = 52;
  ram[2100]  = 255;
  ram[2101]  = 255;
  ram[2102]  = 255;
  ram[2103]  = 255;
  ram[2104]  = 255;
  ram[2105]  = 255;
  ram[2106]  = 255;
  ram[2107]  = 255;
  ram[2108]  = 255;
  ram[2109]  = 255;
  ram[2110]  = 255;
  ram[2111]  = 255;
  ram[2112]  = 255;
  ram[2113]  = 195;
  ram[2114]  = 0;
  ram[2115]  = 0;
  ram[2116]  = 122;
  ram[2117]  = 255;
  ram[2118]  = 255;
  ram[2119]  = 255;
  ram[2120]  = 255;
  ram[2121]  = 255;
  ram[2122]  = 255;
  ram[2123]  = 255;
  ram[2124]  = 255;
  ram[2125]  = 221;
  ram[2126]  = 0;
  ram[2127]  = 0;
  ram[2128]  = 87;
  ram[2129]  = 255;
  ram[2130]  = 255;
  ram[2131]  = 255;
  ram[2132]  = 255;
  ram[2133]  = 71;
  ram[2134]  = 0;
  ram[2135]  = 71;
  ram[2136]  = 255;
  ram[2137]  = 255;
  ram[2138]  = 255;
  ram[2139]  = 255;
  ram[2140]  = 255;
  ram[2141]  = 255;
  ram[2142]  = 255;
  ram[2143]  = 255;
  ram[2144]  = 255;
  ram[2145]  = 255;
  ram[2146]  = 255;
  ram[2147]  = 255;
  ram[2148]  = 255;
  ram[2149]  = 255;
  ram[2150]  = 255;
  ram[2151]  = 255;
  ram[2152]  = 255;
  ram[2153]  = 255;
  ram[2154]  = 255;
  ram[2155]  = 255;
  ram[2156]  = 255;
  ram[2157]  = 255;
  ram[2158]  = 255;
  ram[2159]  = 255;
  ram[2160]  = 255;
  ram[2161]  = 255;
  ram[2162]  = 255;
  ram[2163]  = 255;
  ram[2164]  = 255;
  ram[2165]  = 255;
  ram[2166]  = 255;
  ram[2167]  = 255;
  ram[2168]  = 255;
  ram[2169]  = 255;
  ram[2170]  = 255;
  ram[2171]  = 255;
  ram[2172]  = 255;
  ram[2173]  = 255;
  ram[2174]  = 255;
  ram[2175]  = 255;
  ram[2176]  = 236;
  ram[2177]  = 35;
  ram[2178]  = 0;
  ram[2179]  = 0;
  ram[2180]  = 71;
  ram[2181]  = 236;
  ram[2182]  = 255;
  ram[2183]  = 255;
  ram[2184]  = 255;
  ram[2185]  = 255;
  ram[2186]  = 255;
  ram[2187]  = 255;
  ram[2188]  = 255;
  ram[2189]  = 255;
  ram[2190]  = 236;
  ram[2191]  = 255;
  ram[2192]  = 255;
  ram[2193]  = 105;
  ram[2194]  = 0;
  ram[2195]  = 0;
  ram[2196]  = 208;
  ram[2197]  = 255;
  ram[2198]  = 255;
  ram[2199]  = 255;
  ram[2200]  = 255;
  ram[2201]  = 255;
  ram[2202]  = 255;
  ram[2203]  = 255;
  ram[2204]  = 255;
  ram[2205]  = 255;
  ram[2206]  = 52;
  ram[2207]  = 0;
  ram[2208]  = 0;
  ram[2209]  = 221;
  ram[2210]  = 255;
  ram[2211]  = 255;
  ram[2212]  = 255;
  ram[2213]  = 71;
  ram[2214]  = 0;
  ram[2215]  = 71;
  ram[2216]  = 255;
  ram[2217]  = 255;
  ram[2218]  = 255;
  ram[2219]  = 255;
  ram[2220]  = 255;
  ram[2221]  = 255;
  ram[2222]  = 255;
  ram[2223]  = 255;
  ram[2224]  = 255;
  ram[2225]  = 255;
  ram[2226]  = 255;
  ram[2227]  = 255;
  ram[2228]  = 255;
  ram[2229]  = 255;
  ram[2230]  = 255;
  ram[2231]  = 255;
  ram[2232]  = 255;
  ram[2233]  = 255;
  ram[2234]  = 255;
  ram[2235]  = 255;
  ram[2236]  = 255;
  ram[2237]  = 255;
  ram[2238]  = 255;
  ram[2239]  = 255;
  ram[2240]  = 255;
  ram[2241]  = 255;
  ram[2242]  = 255;
  ram[2243]  = 255;
  ram[2244]  = 255;
  ram[2245]  = 255;
  ram[2246]  = 255;
  ram[2247]  = 255;
  ram[2248]  = 255;
  ram[2249]  = 255;
  ram[2250]  = 255;
  ram[2251]  = 255;
  ram[2252]  = 255;
  ram[2253]  = 255;
  ram[2254]  = 255;
  ram[2255]  = 255;
  ram[2256]  = 255;
  ram[2257]  = 208;
  ram[2258]  = 17;
  ram[2259]  = 0;
  ram[2260]  = 0;
  ram[2261]  = 17;
  ram[2262]  = 137;
  ram[2263]  = 208;
  ram[2264]  = 255;
  ram[2265]  = 255;
  ram[2266]  = 255;
  ram[2267]  = 195;
  ram[2268]  = 152;
  ram[2269]  = 52;
  ram[2270]  = 137;
  ram[2271]  = 255;
  ram[2272]  = 236;
  ram[2273]  = 17;
  ram[2274]  = 0;
  ram[2275]  = 35;
  ram[2276]  = 255;
  ram[2277]  = 255;
  ram[2278]  = 255;
  ram[2279]  = 255;
  ram[2280]  = 255;
  ram[2281]  = 255;
  ram[2282]  = 255;
  ram[2283]  = 255;
  ram[2284]  = 255;
  ram[2285]  = 255;
  ram[2286]  = 167;
  ram[2287]  = 0;
  ram[2288]  = 0;
  ram[2289]  = 137;
  ram[2290]  = 255;
  ram[2291]  = 255;
  ram[2292]  = 255;
  ram[2293]  = 71;
  ram[2294]  = 0;
  ram[2295]  = 71;
  ram[2296]  = 255;
  ram[2297]  = 255;
  ram[2298]  = 255;
  ram[2299]  = 255;
  ram[2300]  = 255;
  ram[2301]  = 255;
  ram[2302]  = 255;
  ram[2303]  = 255;
  ram[2304]  = 255;
  ram[2305]  = 255;
  ram[2306]  = 255;
  ram[2307]  = 255;
  ram[2308]  = 255;
  ram[2309]  = 255;
  ram[2310]  = 255;
  ram[2311]  = 255;
  ram[2312]  = 255;
  ram[2313]  = 255;
  ram[2314]  = 255;
  ram[2315]  = 255;
  ram[2316]  = 255;
  ram[2317]  = 255;
  ram[2318]  = 255;
  ram[2319]  = 255;
  ram[2320]  = 255;
  ram[2321]  = 255;
  ram[2322]  = 255;
  ram[2323]  = 255;
  ram[2324]  = 255;
  ram[2325]  = 255;
  ram[2326]  = 255;
  ram[2327]  = 255;
  ram[2328]  = 255;
  ram[2329]  = 255;
  ram[2330]  = 255;
  ram[2331]  = 255;
  ram[2332]  = 255;
  ram[2333]  = 255;
  ram[2334]  = 255;
  ram[2335]  = 255;
  ram[2336]  = 255;
  ram[2337]  = 255;
  ram[2338]  = 208;
  ram[2339]  = 52;
  ram[2340]  = 0;
  ram[2341]  = 0;
  ram[2342]  = 0;
  ram[2343]  = 0;
  ram[2344]  = 0;
  ram[2345]  = 0;
  ram[2346]  = 0;
  ram[2347]  = 0;
  ram[2348]  = 0;
  ram[2349]  = 0;
  ram[2350]  = 137;
  ram[2351]  = 255;
  ram[2352]  = 167;
  ram[2353]  = 0;
  ram[2354]  = 0;
  ram[2355]  = 137;
  ram[2356]  = 255;
  ram[2357]  = 255;
  ram[2358]  = 255;
  ram[2359]  = 255;
  ram[2360]  = 255;
  ram[2361]  = 255;
  ram[2362]  = 255;
  ram[2363]  = 255;
  ram[2364]  = 255;
  ram[2365]  = 255;
  ram[2366]  = 236;
  ram[2367]  = 0;
  ram[2368]  = 0;
  ram[2369]  = 35;
  ram[2370]  = 255;
  ram[2371]  = 255;
  ram[2372]  = 255;
  ram[2373]  = 71;
  ram[2374]  = 0;
  ram[2375]  = 71;
  ram[2376]  = 255;
  ram[2377]  = 255;
  ram[2378]  = 255;
  ram[2379]  = 255;
  ram[2380]  = 255;
  ram[2381]  = 255;
  ram[2382]  = 255;
  ram[2383]  = 255;
  ram[2384]  = 255;
  ram[2385]  = 255;
  ram[2386]  = 255;
  ram[2387]  = 255;
  ram[2388]  = 255;
  ram[2389]  = 255;
  ram[2390]  = 255;
  ram[2391]  = 255;
  ram[2392]  = 255;
  ram[2393]  = 255;
  ram[2394]  = 255;
  ram[2395]  = 255;
  ram[2396]  = 255;
  ram[2397]  = 255;
  ram[2398]  = 255;
  ram[2399]  = 255;
  ram[2400]  = 255;
  ram[2401]  = 255;
  ram[2402]  = 255;
  ram[2403]  = 255;
  ram[2404]  = 255;
  ram[2405]  = 255;
  ram[2406]  = 255;
  ram[2407]  = 255;
  ram[2408]  = 255;
  ram[2409]  = 255;
  ram[2410]  = 255;
  ram[2411]  = 255;
  ram[2412]  = 255;
  ram[2413]  = 255;
  ram[2414]  = 255;
  ram[2415]  = 255;
  ram[2416]  = 255;
  ram[2417]  = 255;
  ram[2418]  = 255;
  ram[2419]  = 255;
  ram[2420]  = 167;
  ram[2421]  = 52;
  ram[2422]  = 0;
  ram[2423]  = 0;
  ram[2424]  = 0;
  ram[2425]  = 0;
  ram[2426]  = 0;
  ram[2427]  = 0;
  ram[2428]  = 17;
  ram[2429]  = 105;
  ram[2430]  = 208;
  ram[2431]  = 255;
  ram[2432]  = 71;
  ram[2433]  = 0;
  ram[2434]  = 0;
  ram[2435]  = 221;
  ram[2436]  = 255;
  ram[2437]  = 255;
  ram[2438]  = 255;
  ram[2439]  = 255;
  ram[2440]  = 255;
  ram[2441]  = 255;
  ram[2442]  = 255;
  ram[2443]  = 255;
  ram[2444]  = 255;
  ram[2445]  = 255;
  ram[2446]  = 255;
  ram[2447]  = 105;
  ram[2448]  = 0;
  ram[2449]  = 0;
  ram[2450]  = 195;
  ram[2451]  = 255;
  ram[2452]  = 255;
  ram[2453]  = 71;
  ram[2454]  = 0;
  ram[2455]  = 71;
  ram[2456]  = 255;
  ram[2457]  = 255;
  ram[2458]  = 255;
  ram[2459]  = 255;
  ram[2460]  = 255;
  ram[2461]  = 255;
  ram[2462]  = 255;
  ram[2463]  = 255;
  ram[2464]  = 255;
  ram[2465]  = 255;
  ram[2466]  = 255;
  ram[2467]  = 255;
  ram[2468]  = 255;
  ram[2469]  = 255;
  ram[2470]  = 255;
  ram[2471]  = 255;
  ram[2472]  = 255;
  ram[2473]  = 255;
  ram[2474]  = 255;
  ram[2475]  = 255;
  ram[2476]  = 255;
  ram[2477]  = 255;
  ram[2478]  = 255;
  ram[2479]  = 255;
  ram[2480]  = 255;
  ram[2481]  = 255;
  ram[2482]  = 255;
  ram[2483]  = 255;
  ram[2484]  = 255;
  ram[2485]  = 255;
  ram[2486]  = 255;
  ram[2487]  = 255;
  ram[2488]  = 255;
  ram[2489]  = 255;
  ram[2490]  = 255;
  ram[2491]  = 255;
  ram[2492]  = 255;
  ram[2493]  = 255;
  ram[2494]  = 255;
  ram[2495]  = 255;
  ram[2496]  = 255;
  ram[2497]  = 255;
  ram[2498]  = 255;
  ram[2499]  = 255;
  ram[2500]  = 255;
  ram[2501]  = 255;
  ram[2502]  = 236;
  ram[2503]  = 195;
  ram[2504]  = 195;
  ram[2505]  = 195;
  ram[2506]  = 195;
  ram[2507]  = 208;
  ram[2508]  = 255;
  ram[2509]  = 255;
  ram[2510]  = 255;
  ram[2511]  = 255;
  ram[2512]  = 255;
  ram[2513]  = 255;
  ram[2514]  = 255;
  ram[2515]  = 255;
  ram[2516]  = 255;
  ram[2517]  = 255;
  ram[2518]  = 255;
  ram[2519]  = 255;
  ram[2520]  = 255;
  ram[2521]  = 255;
  ram[2522]  = 255;
  ram[2523]  = 255;
  ram[2524]  = 255;
  ram[2525]  = 255;
  ram[2526]  = 255;
  ram[2527]  = 255;
  ram[2528]  = 255;
  ram[2529]  = 255;
  ram[2530]  = 255;
  ram[2531]  = 255;
  ram[2532]  = 255;
  ram[2533]  = 255;
  ram[2534]  = 255;
  ram[2535]  = 255;
  ram[2536]  = 255;
  ram[2537]  = 255;
  ram[2538]  = 255;
  ram[2539]  = 255;
  ram[2540]  = 255;
  ram[2541]  = 255;
  ram[2542]  = 255;
  ram[2543]  = 255;
  ram[2544]  = 255;
  ram[2545]  = 255;
  ram[2546]  = 255;
  ram[2547]  = 255;
  ram[2548]  = 255;
  ram[2549]  = 255;
  ram[2550]  = 255;
  ram[2551]  = 255;
  ram[2552]  = 255;
  ram[2553]  = 255;
  ram[2554]  = 255;
  ram[2555]  = 255;
  ram[2556]  = 255;
  ram[2557]  = 255;
  ram[2558]  = 255;
  ram[2559]  = 255;
  ram[2560]  = 255;
  ram[2561]  = 255;
  ram[2562]  = 255;
  ram[2563]  = 255;
  ram[2564]  = 255;
  ram[2565]  = 255;
  ram[2566]  = 255;
  ram[2567]  = 255;
  ram[2568]  = 255;
  ram[2569]  = 255;
  ram[2570]  = 255;
  ram[2571]  = 255;
  ram[2572]  = 255;
  ram[2573]  = 255;
  ram[2574]  = 255;
  ram[2575]  = 255;
  ram[2576]  = 255;
  ram[2577]  = 255;
  ram[2578]  = 255;
  ram[2579]  = 255;
  ram[2580]  = 255;
  ram[2581]  = 255;
  ram[2582]  = 255;
  ram[2583]  = 255;
  ram[2584]  = 255;
  ram[2585]  = 255;
  ram[2586]  = 255;
  ram[2587]  = 255;
  ram[2588]  = 255;
  ram[2589]  = 255;
  ram[2590]  = 255;
  ram[2591]  = 255;
  ram[2592]  = 255;
  ram[2593]  = 255;
  ram[2594]  = 255;
  ram[2595]  = 255;
  ram[2596]  = 255;
  ram[2597]  = 255;
  ram[2598]  = 255;
  ram[2599]  = 255;
  ram[2600]  = 255;
  ram[2601]  = 255;
  ram[2602]  = 255;
  ram[2603]  = 255;
  ram[2604]  = 255;
  ram[2605]  = 255;
  ram[2606]  = 255;
  ram[2607]  = 255;
  ram[2608]  = 255;
  ram[2609]  = 255;
  ram[2610]  = 255;
  ram[2611]  = 255;
  ram[2612]  = 255;
  ram[2613]  = 255;
  ram[2614]  = 255;
  ram[2615]  = 255;
  ram[2616]  = 255;
  ram[2617]  = 255;
  ram[2618]  = 255;
  ram[2619]  = 255;
  ram[2620]  = 255;
  ram[2621]  = 255;
  ram[2622]  = 255;
  ram[2623]  = 255;
  ram[2624]  = 255;
  ram[2625]  = 255;
  ram[2626]  = 255;
  ram[2627]  = 255;
  ram[2628]  = 255;
  ram[2629]  = 255;
  ram[2630]  = 255;
  ram[2631]  = 255;
  ram[2632]  = 255;
  ram[2633]  = 255;
  ram[2634]  = 255;
  ram[2635]  = 255;
  ram[2636]  = 255;
  ram[2637]  = 255;
  ram[2638]  = 255;
  ram[2639]  = 255;
  ram[2640]  = 255;
  ram[2641]  = 255;
  ram[2642]  = 255;
  ram[2643]  = 255;
  ram[2644]  = 255;
  ram[2645]  = 255;
  ram[2646]  = 255;
  ram[2647]  = 255;
  ram[2648]  = 255;
  ram[2649]  = 255;
  ram[2650]  = 255;
  ram[2651]  = 255;
  ram[2652]  = 255;
  ram[2653]  = 255;
  ram[2654]  = 255;
  ram[2655]  = 255;
  ram[2656]  = 255;
  ram[2657]  = 255;
  ram[2658]  = 255;
  ram[2659]  = 255;
  ram[2660]  = 255;
  ram[2661]  = 255;
  ram[2662]  = 255;
  ram[2663]  = 255;
  ram[2664]  = 255;
  ram[2665]  = 255;
  ram[2666]  = 255;
  ram[2667]  = 255;
  ram[2668]  = 255;
  ram[2669]  = 255;
  ram[2670]  = 255;
  ram[2671]  = 255;
  ram[2672]  = 255;
  ram[2673]  = 255;
  ram[2674]  = 255;
  ram[2675]  = 255;
  ram[2676]  = 255;
  ram[2677]  = 255;
  ram[2678]  = 255;
  ram[2679]  = 255;
  ram[2680]  = 255;
  ram[2681]  = 255;
  ram[2682]  = 255;
  ram[2683]  = 255;
  ram[2684]  = 255;
  ram[2685]  = 255;
  ram[2686]  = 255;
  ram[2687]  = 255;
  ram[2688]  = 255;
  ram[2689]  = 255;
  ram[2690]  = 255;
  ram[2691]  = 255;
  ram[2692]  = 255;
  ram[2693]  = 255;
  ram[2694]  = 255;
  ram[2695]  = 255;
  ram[2696]  = 255;
  ram[2697]  = 255;
  ram[2698]  = 255;
  ram[2699]  = 255;
  ram[2700]  = 255;
  ram[2701]  = 255;
  ram[2702]  = 255;
  ram[2703]  = 255;
  ram[2704]  = 255;
  ram[2705]  = 255;
  ram[2706]  = 255;
  ram[2707]  = 255;
  ram[2708]  = 255;
  ram[2709]  = 255;
  ram[2710]  = 255;
  ram[2711]  = 255;
  ram[2712]  = 255;
  ram[2713]  = 255;
  ram[2714]  = 255;
  ram[2715]  = 255;
  ram[2716]  = 255;
  ram[2717]  = 255;
  ram[2718]  = 255;
  ram[2719]  = 255;
  ram[2720]  = 255;
  ram[2721]  = 255;
  ram[2722]  = 255;
  ram[2723]  = 255;
  ram[2724]  = 255;
  ram[2725]  = 255;
  ram[2726]  = 255;
  ram[2727]  = 255;
  ram[2728]  = 255;
  ram[2729]  = 255;
  ram[2730]  = 255;
  ram[2731]  = 255;
  ram[2732]  = 255;
  ram[2733]  = 255;
  ram[2734]  = 255;
  ram[2735]  = 255;
  ram[2736]  = 255;
  ram[2737]  = 255;
  ram[2738]  = 255;
  ram[2739]  = 255;
  ram[2740]  = 255;
  ram[2741]  = 255;
  ram[2742]  = 255;
  ram[2743]  = 255;
  ram[2744]  = 255;
  ram[2745]  = 255;
  ram[2746]  = 255;
  ram[2747]  = 255;
  ram[2748]  = 255;
  ram[2749]  = 255;
  ram[2750]  = 255;
  ram[2751]  = 255;
  ram[2752]  = 255;
  ram[2753]  = 255;
  ram[2754]  = 255;
  ram[2755]  = 255;
  ram[2756]  = 255;
  ram[2757]  = 255;
  ram[2758]  = 255;
  ram[2759]  = 255;
  ram[2760]  = 255;
  ram[2761]  = 255;
  ram[2762]  = 255;
  ram[2763]  = 255;
  ram[2764]  = 255;
  ram[2765]  = 255;
  ram[2766]  = 255;
  ram[2767]  = 255;
  ram[2768]  = 255;
  ram[2769]  = 255;
  ram[2770]  = 255;
  ram[2771]  = 255;
  ram[2772]  = 255;
  ram[2773]  = 255;
  ram[2774]  = 255;
  ram[2775]  = 255;
  ram[2776]  = 255;
  ram[2777]  = 255;
  ram[2778]  = 255;
  ram[2779]  = 255;
  ram[2780]  = 255;
  ram[2781]  = 255;
  ram[2782]  = 255;
  ram[2783]  = 255;
  ram[2784]  = 255;
  ram[2785]  = 255;
  ram[2786]  = 255;
  ram[2787]  = 255;
  ram[2788]  = 255;
  ram[2789]  = 255;
  ram[2790]  = 255;
  ram[2791]  = 255;
  ram[2792]  = 255;
  ram[2793]  = 255;
  ram[2794]  = 255;
  ram[2795]  = 255;
  ram[2796]  = 255;
  ram[2797]  = 255;
  ram[2798]  = 255;
  ram[2799]  = 255;
  ram[2800]  = 255;
  ram[2801]  = 255;
  ram[2802]  = 255;
  ram[2803]  = 255;
  ram[2804]  = 255;
  ram[2805]  = 255;
  ram[2806]  = 255;
  ram[2807]  = 255;
  ram[2808]  = 255;
  ram[2809]  = 255;
  ram[2810]  = 255;
  ram[2811]  = 255;
  ram[2812]  = 255;
  ram[2813]  = 255;
  ram[2814]  = 255;
  ram[2815]  = 255;
  ram[2816]  = 255;
  ram[2817]  = 255;
  ram[2818]  = 255;
  ram[2819]  = 255;
  ram[2820]  = 255;
  ram[2821]  = 255;
  ram[2822]  = 255;
  ram[2823]  = 255;
  ram[2824]  = 255;
  ram[2825]  = 255;
  ram[2826]  = 255;
  ram[2827]  = 255;
  ram[2828]  = 255;
  ram[2829]  = 255;
  ram[2830]  = 255;
  ram[2831]  = 255;
  ram[2832]  = 255;
  ram[2833]  = 255;
  ram[2834]  = 255;
  ram[2835]  = 255;
  ram[2836]  = 255;
  ram[2837]  = 255;
  ram[2838]  = 255;
  ram[2839]  = 255;
  ram[2840]  = 255;
  ram[2841]  = 255;
  ram[2842]  = 255;
  ram[2843]  = 255;
  ram[2844]  = 255;
  ram[2845]  = 255;
  ram[2846]  = 255;
  ram[2847]  = 255;
  ram[2848]  = 255;
  ram[2849]  = 255;
  ram[2850]  = 255;
  ram[2851]  = 255;
  ram[2852]  = 255;
  ram[2853]  = 255;
  ram[2854]  = 255;
  ram[2855]  = 255;
  ram[2856]  = 255;
  ram[2857]  = 255;
  ram[2858]  = 255;
  ram[2859]  = 255;
  ram[2860]  = 255;
  ram[2861]  = 255;
  ram[2862]  = 255;
  ram[2863]  = 255;
  ram[2864]  = 255;
  ram[2865]  = 255;
  ram[2866]  = 255;
  ram[2867]  = 255;
  ram[2868]  = 255;
  ram[2869]  = 255;
  ram[2870]  = 255;
  ram[2871]  = 255;
  ram[2872]  = 255;
  ram[2873]  = 255;
  ram[2874]  = 255;
  ram[2875]  = 255;
  ram[2876]  = 255;
  ram[2877]  = 255;
  ram[2878]  = 255;
  ram[2879]  = 255;
  ram[2880]  = 255;
  ram[2881]  = 255;
  ram[2882]  = 255;
  ram[2883]  = 255;
  ram[2884]  = 255;
  ram[2885]  = 255;
  ram[2886]  = 255;
  ram[2887]  = 255;
  ram[2888]  = 255;
  ram[2889]  = 255;
  ram[2890]  = 255;
  ram[2891]  = 255;
  ram[2892]  = 255;
  ram[2893]  = 255;
  ram[2894]  = 255;
  ram[2895]  = 255;
  ram[2896]  = 255;
  ram[2897]  = 255;
  ram[2898]  = 255;
  ram[2899]  = 255;
  ram[2900]  = 255;
  ram[2901]  = 255;
  ram[2902]  = 255;
  ram[2903]  = 255;
  ram[2904]  = 255;
  ram[2905]  = 255;
  ram[2906]  = 255;
  ram[2907]  = 255;
  ram[2908]  = 255;
  ram[2909]  = 255;
  ram[2910]  = 255;
  ram[2911]  = 255;
  ram[2912]  = 255;
  ram[2913]  = 255;
  ram[2914]  = 255;
  ram[2915]  = 255;
  ram[2916]  = 255;
  ram[2917]  = 255;
  ram[2918]  = 255;
  ram[2919]  = 255;
  ram[2920]  = 255;
  ram[2921]  = 255;
  ram[2922]  = 255;
  ram[2923]  = 255;
  ram[2924]  = 255;
  ram[2925]  = 255;
  ram[2926]  = 255;
  ram[2927]  = 255;
  ram[2928]  = 255;
  ram[2929]  = 255;
  ram[2930]  = 255;
  ram[2931]  = 255;
  ram[2932]  = 255;
  ram[2933]  = 255;
  ram[2934]  = 255;
  ram[2935]  = 255;
  ram[2936]  = 255;
  ram[2937]  = 255;
  ram[2938]  = 255;
  ram[2939]  = 255;
  ram[2940]  = 255;
  ram[2941]  = 255;
  ram[2942]  = 255;
  ram[2943]  = 255;
  ram[2944]  = 255;
  ram[2945]  = 255;
  ram[2946]  = 255;
  ram[2947]  = 255;
  ram[2948]  = 255;
  ram[2949]  = 255;
  ram[2950]  = 255;
  ram[2951]  = 255;
  ram[2952]  = 255;
  ram[2953]  = 255;
  ram[2954]  = 255;
  ram[2955]  = 255;
  ram[2956]  = 255;
  ram[2957]  = 255;
  ram[2958]  = 255;
  ram[2959]  = 255;
  ram[2960]  = 255;
  ram[2961]  = 255;
  ram[2962]  = 255;
  ram[2963]  = 255;
  ram[2964]  = 255;
  ram[2965]  = 255;
  ram[2966]  = 255;
  ram[2967]  = 255;
  ram[2968]  = 255;
  ram[2969]  = 255;
  ram[2970]  = 255;
  ram[2971]  = 255;
  ram[2972]  = 255;
  ram[2973]  = 255;
  ram[2974]  = 255;
  ram[2975]  = 255;
  ram[2976]  = 255;
  ram[2977]  = 255;
  ram[2978]  = 255;
  ram[2979]  = 255;
  ram[2980]  = 255;
  ram[2981]  = 255;
  ram[2982]  = 255;
  ram[2983]  = 255;
  ram[2984]  = 255;
  ram[2985]  = 255;
  ram[2986]  = 255;
  ram[2987]  = 255;
  ram[2988]  = 255;
  ram[2989]  = 255;
  ram[2990]  = 255;
  ram[2991]  = 255;
  ram[2992]  = 255;
  ram[2993]  = 255;
  ram[2994]  = 255;
  ram[2995]  = 255;
  ram[2996]  = 255;
  ram[2997]  = 255;
  ram[2998]  = 255;
  ram[2999]  = 255;
  ram[3000]  = 255;
  ram[3001]  = 255;
  ram[3002]  = 255;
  ram[3003]  = 255;
  ram[3004]  = 255;
  ram[3005]  = 255;
  ram[3006]  = 255;
  ram[3007]  = 255;
  ram[3008]  = 255;
  ram[3009]  = 255;
  ram[3010]  = 255;
  ram[3011]  = 255;
  ram[3012]  = 255;
  ram[3013]  = 255;
  ram[3014]  = 255;
  ram[3015]  = 255;
  ram[3016]  = 255;
  ram[3017]  = 255;
  ram[3018]  = 255;
  ram[3019]  = 255;
  ram[3020]  = 255;
  ram[3021]  = 255;
  ram[3022]  = 255;
  ram[3023]  = 255;
  ram[3024]  = 255;
  ram[3025]  = 255;
  ram[3026]  = 255;
  ram[3027]  = 255;
  ram[3028]  = 255;
  ram[3029]  = 255;
  ram[3030]  = 255;
  ram[3031]  = 255;
  ram[3032]  = 255;
  ram[3033]  = 255;
  ram[3034]  = 255;
  ram[3035]  = 255;
  ram[3036]  = 255;
  ram[3037]  = 255;
  ram[3038]  = 255;
  ram[3039]  = 255;
  ram[3040]  = 255;
  ram[3041]  = 255;
  ram[3042]  = 255;
  ram[3043]  = 255;
  ram[3044]  = 255;
  ram[3045]  = 255;
  ram[3046]  = 255;
  ram[3047]  = 255;
  ram[3048]  = 255;
  ram[3049]  = 255;
  ram[3050]  = 255;
  ram[3051]  = 255;
  ram[3052]  = 255;
  ram[3053]  = 255;
  ram[3054]  = 255;
  ram[3055]  = 255;
  ram[3056]  = 255;
  ram[3057]  = 255;
  ram[3058]  = 255;
  ram[3059]  = 255;
  ram[3060]  = 255;
  ram[3061]  = 255;
  ram[3062]  = 255;
  ram[3063]  = 255;
  ram[3064]  = 255;
  ram[3065]  = 255;
  ram[3066]  = 255;
  ram[3067]  = 255;
  ram[3068]  = 255;
  ram[3069]  = 255;
  ram[3070]  = 255;
  ram[3071]  = 255;
  ram[3072]  = 255;
  ram[3073]  = 255;
  ram[3074]  = 255;
  ram[3075]  = 255;
  ram[3076]  = 255;
  ram[3077]  = 255;
  ram[3078]  = 255;
  ram[3079]  = 255;
  ram[3080]  = 255;
  ram[3081]  = 255;
  ram[3082]  = 255;
  ram[3083]  = 255;
  ram[3084]  = 255;
  ram[3085]  = 255;
  ram[3086]  = 255;
  ram[3087]  = 255;
  ram[3088]  = 255;
  ram[3089]  = 255;
  ram[3090]  = 255;
  ram[3091]  = 255;
  ram[3092]  = 255;
  ram[3093]  = 255;
  ram[3094]  = 255;
  ram[3095]  = 255;
  ram[3096]  = 255;
  ram[3097]  = 255;
  ram[3098]  = 255;
  ram[3099]  = 255;
  ram[3100]  = 255;
  ram[3101]  = 255;
  ram[3102]  = 255;
  ram[3103]  = 255;
  ram[3104]  = 255;
  ram[3105]  = 255;
  ram[3106]  = 255;
  ram[3107]  = 255;
  ram[3108]  = 255;
  ram[3109]  = 255;
  ram[3110]  = 255;
  ram[3111]  = 255;
  ram[3112]  = 255;
  ram[3113]  = 255;
  ram[3114]  = 255;
  ram[3115]  = 255;
  ram[3116]  = 255;
  ram[3117]  = 255;
  ram[3118]  = 255;
  ram[3119]  = 255;
  ram[3120]  = 255;
  ram[3121]  = 255;
  ram[3122]  = 255;
  ram[3123]  = 255;
  ram[3124]  = 255;
  ram[3125]  = 255;
  ram[3126]  = 255;
  ram[3127]  = 255;
  ram[3128]  = 255;
  ram[3129]  = 255;
  ram[3130]  = 255;
  ram[3131]  = 255;
  ram[3132]  = 255;
  ram[3133]  = 255;
  ram[3134]  = 255;
  ram[3135]  = 255;
  ram[3136]  = 255;
  ram[3137]  = 255;
  ram[3138]  = 255;
  ram[3139]  = 255;
  ram[3140]  = 255;
  ram[3141]  = 255;
  ram[3142]  = 255;
  ram[3143]  = 255;
  ram[3144]  = 255;
  ram[3145]  = 255;
  ram[3146]  = 255;
  ram[3147]  = 255;
  ram[3148]  = 255;
  ram[3149]  = 255;
  ram[3150]  = 255;
  ram[3151]  = 255;
  ram[3152]  = 255;
  ram[3153]  = 255;
  ram[3154]  = 255;
  ram[3155]  = 255;
  ram[3156]  = 255;
  ram[3157]  = 255;
  ram[3158]  = 255;
  ram[3159]  = 255;
  ram[3160]  = 255;
  ram[3161]  = 255;
  ram[3162]  = 255;
  ram[3163]  = 255;
  ram[3164]  = 255;
  ram[3165]  = 255;
  ram[3166]  = 255;
  ram[3167]  = 255;
  ram[3168]  = 255;
  ram[3169]  = 255;
  ram[3170]  = 255;
  ram[3171]  = 255;
  ram[3172]  = 255;
  ram[3173]  = 255;
  ram[3174]  = 255;
  ram[3175]  = 255;
  ram[3176]  = 255;
  ram[3177]  = 255;
  ram[3178]  = 255;
  ram[3179]  = 255;
  ram[3180]  = 255;
  ram[3181]  = 255;
  ram[3182]  = 255;
  ram[3183]  = 255;
  ram[3184]  = 255;
  ram[3185]  = 255;
  ram[3186]  = 255;
  ram[3187]  = 255;
  ram[3188]  = 255;
  ram[3189]  = 255;
  ram[3190]  = 255;
  ram[3191]  = 255;
  ram[3192]  = 255;
  ram[3193]  = 255;
  ram[3194]  = 255;
  ram[3195]  = 255;
  ram[3196]  = 255;
  ram[3197]  = 255;
  ram[3198]  = 255;
  ram[3199]  = 255;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
