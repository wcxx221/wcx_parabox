module rom_dist_b(clock, address, q);       // ROM-stored RGB bitmap for level destination
input clock;
output [7:0] q;
input [8:0] address;
reg [7:0] dout;
reg [7:0] ram [511:0];
assign q = dout;

initial begin
  ram[0]  = 255;
  ram[1]  = 255;
  ram[2]  = 255;
  ram[3]  = 255;
  ram[4]  = 255;
  ram[5]  = 255;
  ram[6]  = 255;
  ram[7]  = 0;
  ram[8]  = 0;
  ram[9]  = 0;
  ram[10]  = 0;
  ram[11]  = 0;
  ram[12]  = 255;
  ram[13]  = 255;
  ram[14]  = 255;
  ram[15]  = 255;
  ram[16]  = 255;
  ram[17]  = 255;
  ram[18]  = 255;
  ram[19]  = 255;
  ram[20]  = 255;
  ram[21]  = 255;
  ram[22]  = 255;
  ram[23]  = 255;
  ram[24]  = 255;
  ram[25]  = 0;
  ram[26]  = 0;
  ram[27]  = 0;
  ram[28]  = 0;
  ram[29]  = 0;
  ram[30]  = 0;
  ram[31]  = 0;
  ram[32]  = 0;
  ram[33]  = 0;
  ram[34]  = 255;
  ram[35]  = 255;
  ram[36]  = 255;
  ram[37]  = 255;
  ram[38]  = 255;
  ram[39]  = 255;
  ram[40]  = 255;
  ram[41]  = 255;
  ram[42]  = 255;
  ram[43]  = 0;
  ram[44]  = 0;
  ram[45]  = 0;
  ram[46]  = 0;
  ram[47]  = 0;
  ram[48]  = 0;
  ram[49]  = 0;
  ram[50]  = 0;
  ram[51]  = 0;
  ram[52]  = 0;
  ram[53]  = 0;
  ram[54]  = 0;
  ram[55]  = 0;
  ram[56]  = 255;
  ram[57]  = 255;
  ram[58]  = 255;
  ram[59]  = 255;
  ram[60]  = 255;
  ram[61]  = 255;
  ram[62]  = 0;
  ram[63]  = 0;
  ram[64]  = 0;
  ram[65]  = 0;
  ram[66]  = 0;
  ram[67]  = 0;
  ram[68]  = 0;
  ram[69]  = 0;
  ram[70]  = 0;
  ram[71]  = 0;
  ram[72]  = 0;
  ram[73]  = 0;
  ram[74]  = 0;
  ram[75]  = 0;
  ram[76]  = 0;
  ram[77]  = 255;
  ram[78]  = 255;
  ram[79]  = 255;
  ram[80]  = 255;
  ram[81]  = 255;
  ram[82]  = 0;
  ram[83]  = 0;
  ram[84]  = 0;
  ram[85]  = 0;
  ram[86]  = 0;
  ram[87]  = 0;
  ram[88]  = 0;
  ram[89]  = 0;
  ram[90]  = 0;
  ram[91]  = 0;
  ram[92]  = 0;
  ram[93]  = 0;
  ram[94]  = 0;
  ram[95]  = 0;
  ram[96]  = 0;
  ram[97]  = 255;
  ram[98]  = 255;
  ram[99]  = 255;
  ram[100]  = 255;
  ram[101]  = 0;
  ram[102]  = 0;
  ram[103]  = 0;
  ram[104]  = 0;
  ram[105]  = 0;
  ram[106]  = 0;
  ram[107]  = 0;
  ram[108]  = 255;
  ram[109]  = 255;
  ram[110]  = 255;
  ram[111]  = 0;
  ram[112]  = 0;
  ram[113]  = 0;
  ram[114]  = 0;
  ram[115]  = 0;
  ram[116]  = 0;
  ram[117]  = 0;
  ram[118]  = 255;
  ram[119]  = 255;
  ram[120]  = 255;
  ram[121]  = 0;
  ram[122]  = 0;
  ram[123]  = 0;
  ram[124]  = 0;
  ram[125]  = 0;
  ram[126]  = 255;
  ram[127]  = 255;
  ram[128]  = 255;
  ram[129]  = 255;
  ram[130]  = 255;
  ram[131]  = 255;
  ram[132]  = 255;
  ram[133]  = 0;
  ram[134]  = 0;
  ram[135]  = 0;
  ram[136]  = 0;
  ram[137]  = 0;
  ram[138]  = 255;
  ram[139]  = 255;
  ram[140]  = 0;
  ram[141]  = 0;
  ram[142]  = 0;
  ram[143]  = 0;
  ram[144]  = 0;
  ram[145]  = 0;
  ram[146]  = 255;
  ram[147]  = 255;
  ram[148]  = 255;
  ram[149]  = 255;
  ram[150]  = 255;
  ram[151]  = 255;
  ram[152]  = 255;
  ram[153]  = 0;
  ram[154]  = 0;
  ram[155]  = 0;
  ram[156]  = 0;
  ram[157]  = 0;
  ram[158]  = 0;
  ram[159]  = 255;
  ram[160]  = 0;
  ram[161]  = 0;
  ram[162]  = 0;
  ram[163]  = 0;
  ram[164]  = 0;
  ram[165]  = 255;
  ram[166]  = 255;
  ram[167]  = 255;
  ram[168]  = 255;
  ram[169]  = 255;
  ram[170]  = 255;
  ram[171]  = 255;
  ram[172]  = 255;
  ram[173]  = 255;
  ram[174]  = 0;
  ram[175]  = 0;
  ram[176]  = 0;
  ram[177]  = 0;
  ram[178]  = 0;
  ram[179]  = 255;
  ram[180]  = 0;
  ram[181]  = 0;
  ram[182]  = 0;
  ram[183]  = 0;
  ram[184]  = 0;
  ram[185]  = 255;
  ram[186]  = 255;
  ram[187]  = 255;
  ram[188]  = 255;
  ram[189]  = 255;
  ram[190]  = 255;
  ram[191]  = 255;
  ram[192]  = 255;
  ram[193]  = 255;
  ram[194]  = 0;
  ram[195]  = 0;
  ram[196]  = 0;
  ram[197]  = 0;
  ram[198]  = 0;
  ram[199]  = 255;
  ram[200]  = 0;
  ram[201]  = 0;
  ram[202]  = 0;
  ram[203]  = 0;
  ram[204]  = 0;
  ram[205]  = 255;
  ram[206]  = 255;
  ram[207]  = 255;
  ram[208]  = 255;
  ram[209]  = 255;
  ram[210]  = 255;
  ram[211]  = 255;
  ram[212]  = 255;
  ram[213]  = 255;
  ram[214]  = 0;
  ram[215]  = 0;
  ram[216]  = 0;
  ram[217]  = 0;
  ram[218]  = 0;
  ram[219]  = 255;
  ram[220]  = 0;
  ram[221]  = 0;
  ram[222]  = 0;
  ram[223]  = 0;
  ram[224]  = 0;
  ram[225]  = 255;
  ram[226]  = 255;
  ram[227]  = 255;
  ram[228]  = 255;
  ram[229]  = 255;
  ram[230]  = 255;
  ram[231]  = 255;
  ram[232]  = 255;
  ram[233]  = 255;
  ram[234]  = 0;
  ram[235]  = 0;
  ram[236]  = 0;
  ram[237]  = 0;
  ram[238]  = 0;
  ram[239]  = 255;
  ram[240]  = 0;
  ram[241]  = 0;
  ram[242]  = 0;
  ram[243]  = 0;
  ram[244]  = 0;
  ram[245]  = 0;
  ram[246]  = 255;
  ram[247]  = 255;
  ram[248]  = 255;
  ram[249]  = 255;
  ram[250]  = 255;
  ram[251]  = 255;
  ram[252]  = 255;
  ram[253]  = 0;
  ram[254]  = 0;
  ram[255]  = 0;
  ram[256]  = 0;
  ram[257]  = 0;
  ram[258]  = 0;
  ram[259]  = 255;
  ram[260]  = 255;
  ram[261]  = 0;
  ram[262]  = 0;
  ram[263]  = 0;
  ram[264]  = 0;
  ram[265]  = 0;
  ram[266]  = 255;
  ram[267]  = 255;
  ram[268]  = 255;
  ram[269]  = 255;
  ram[270]  = 255;
  ram[271]  = 255;
  ram[272]  = 255;
  ram[273]  = 0;
  ram[274]  = 0;
  ram[275]  = 0;
  ram[276]  = 0;
  ram[277]  = 0;
  ram[278]  = 255;
  ram[279]  = 255;
  ram[280]  = 255;
  ram[281]  = 0;
  ram[282]  = 0;
  ram[283]  = 0;
  ram[284]  = 0;
  ram[285]  = 0;
  ram[286]  = 0;
  ram[287]  = 0;
  ram[288]  = 255;
  ram[289]  = 255;
  ram[290]  = 255;
  ram[291]  = 0;
  ram[292]  = 0;
  ram[293]  = 0;
  ram[294]  = 0;
  ram[295]  = 0;
  ram[296]  = 0;
  ram[297]  = 0;
  ram[298]  = 255;
  ram[299]  = 255;
  ram[300]  = 255;
  ram[301]  = 255;
  ram[302]  = 0;
  ram[303]  = 0;
  ram[304]  = 0;
  ram[305]  = 0;
  ram[306]  = 0;
  ram[307]  = 0;
  ram[308]  = 0;
  ram[309]  = 0;
  ram[310]  = 0;
  ram[311]  = 0;
  ram[312]  = 0;
  ram[313]  = 0;
  ram[314]  = 0;
  ram[315]  = 0;
  ram[316]  = 0;
  ram[317]  = 255;
  ram[318]  = 255;
  ram[319]  = 255;
  ram[320]  = 255;
  ram[321]  = 255;
  ram[322]  = 0;
  ram[323]  = 0;
  ram[324]  = 0;
  ram[325]  = 0;
  ram[326]  = 0;
  ram[327]  = 0;
  ram[328]  = 0;
  ram[329]  = 0;
  ram[330]  = 0;
  ram[331]  = 0;
  ram[332]  = 0;
  ram[333]  = 0;
  ram[334]  = 0;
  ram[335]  = 0;
  ram[336]  = 0;
  ram[337]  = 255;
  ram[338]  = 255;
  ram[339]  = 255;
  ram[340]  = 255;
  ram[341]  = 255;
  ram[342]  = 255;
  ram[343]  = 0;
  ram[344]  = 0;
  ram[345]  = 0;
  ram[346]  = 0;
  ram[347]  = 0;
  ram[348]  = 0;
  ram[349]  = 0;
  ram[350]  = 0;
  ram[351]  = 0;
  ram[352]  = 0;
  ram[353]  = 0;
  ram[354]  = 0;
  ram[355]  = 0;
  ram[356]  = 255;
  ram[357]  = 255;
  ram[358]  = 255;
  ram[359]  = 255;
  ram[360]  = 255;
  ram[361]  = 255;
  ram[362]  = 255;
  ram[363]  = 255;
  ram[364]  = 255;
  ram[365]  = 0;
  ram[366]  = 0;
  ram[367]  = 0;
  ram[368]  = 0;
  ram[369]  = 0;
  ram[370]  = 0;
  ram[371]  = 0;
  ram[372]  = 0;
  ram[373]  = 0;
  ram[374]  = 255;
  ram[375]  = 255;
  ram[376]  = 255;
  ram[377]  = 255;
  ram[378]  = 255;
  ram[379]  = 255;
  ram[380]  = 255;
  ram[381]  = 255;
  ram[382]  = 255;
  ram[383]  = 255;
  ram[384]  = 255;
  ram[385]  = 255;
  ram[386]  = 255;
  ram[387]  = 0;
  ram[388]  = 0;
  ram[389]  = 0;
  ram[390]  = 0;
  ram[391]  = 0;
  ram[392]  = 255;
  ram[393]  = 255;
  ram[394]  = 255;
  ram[395]  = 255;
  ram[396]  = 255;
  ram[397]  = 255;
  ram[398]  = 255;
  ram[399]  = 255;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
